module ctrl_blk_2(
	input 		fifo_empty,
	input 		clk_2,
	input 		reset_n,
	output reg 	zero_sel,
	output reg 	rd_fifo,
	output reg 	ram_ena,
	output reg 	ram_wr_n
	);


enum reg {
read_idle = 1'b0,
read = 1'b1,
read_xx	= 'x
} read_ps, read_ns;

enum reg [1:0] {
ram_write_idle = 2'b00,
ram_write = 2'b01,
ram_write_wait = 2'b10,
ram_write_xx = 'x
} ram_write_ps, ram_write_ns;

enum reg [2:0] {idle		= 3'b000,
		byte_0		= 3'b001,
          	byte_1		= 3'b010,
          	byte_2		= 3'b011,
          	byte_3		= 3'b100,
          	byte_xx	= 'x} byte_cnt_ps, byte_cnt_ns;



//************************************************************
//sm #1 read fifo active or not  
//************************************************************
always_ff @(posedge clk_2, negedge reset_n)
    	if (!reset_n) read_ps <= read_idle;        //after reset, go to state 'not_complete'
    	else          read_ps <= read_ns;        //else, go to next state

always_comb begin
    	read_ns = read_xx;   //default assignments;
	rd_fifo = 1'b0;
    	unique case (read_ps)
     		read_idle:
			if (!fifo_empty)  read_ns = read;
			else read_ns = read_idle;
     		read:
			begin
				rd_fifo = 1'b1;	
				read_ns = read_idle;
			end
    	endcase
end//always_comb


always_comb begin
	if (byte_cnt_ps == byte_0)		
		zero_sel = 1'b1;
	else 
		zero_sel = 1'b0;
end

//************************************************************
//sm #2  Is it the first byte?
//************************************************************
//always_ff @(posedge clk_2, negedge reset_n)
 //   	if (!reset_n) first_byte_ps <= first_byte_n;        //after reset, go to state 'first_byte_n'
 //   	else          first_byte_ps <= first_byte_ns;        //else, go to next state

//always_comb begin
//    	first_byte_ns = first_byte_xx;   //default assignments;
//	zero_sel = 1'b0;
//    	unique case (first_byte_ps)
 //    		first_byte_n:
//			if (byte_cnt_ns == byte_1) first_byte_ns = first_byte;
//			else first_byte_ns = first_byte_n;
//     		first_byte:  
//			begin
//				first_byte_ns = first_byte_n;
//				zero_sel = 1'b1;
//			end
//    	endcase
//end

//************************************************************
//sm #3  what byte
//************************************************************
always_ff @(posedge clk_2, negedge reset_n)
    	if (!reset_n) byte_cnt_ps <= byte_0;        //after reset, go to state 'not_complete'
    	else          byte_cnt_ps <= byte_cnt_ns;   //else, go to next state

always_comb begin
    	byte_cnt_ns = byte_xx;   //default assignments; 
    	case (byte_cnt_ps)
     		byte_0:
			if (read_ps == read & (!fifo_empty)) byte_cnt_ns = byte_1;
			else byte_cnt_ns = byte_0;
     		byte_1:
			if (read_ps == read & (!fifo_empty)) byte_cnt_ns = byte_2;
			else byte_cnt_ns = byte_1;
     		byte_2:
			if (read_ps == read & (!fifo_empty)) byte_cnt_ns = byte_3;
			else byte_cnt_ns = byte_2;
     		byte_3:
			if (read_ps == read & (!fifo_empty)) byte_cnt_ns = byte_0;
			else byte_cnt_ns = byte_3;
    	endcase
end



//************************************************************
//sm #4  write to ram?
//************************************************************
always_ff @(posedge clk_2, negedge reset_n)
    	if (!reset_n) ram_write_ps <= ram_write_idle;  	//after reset, go to state 'first_byte_n'
    	else          ram_write_ps <= ram_write_ns;   	//else, go to next state

always_comb begin
    	ram_write_ns = ram_write_xx;   //default assignments;
	ram_ena = 1'b0;
	ram_wr_n = 1'b1;
    	case (ram_write_ps)

     		ram_write_idle:
			if ((byte_cnt_ps == byte_3) && (read_ps == read))  ram_write_ns = ram_write;
			else ram_write_ns = ram_write_idle;
     		ram_write:
			begin
				ram_write_ns = ram_write_wait;
				ram_wr_n = 1'b0;
			end
     		ram_write_wait:
			begin
				ram_write_ns = ram_write_idle;
				ram_ena = 1'b1;
			end
    	endcase
end//always

endmodule
