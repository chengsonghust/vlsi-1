
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, n14, n15, n16, n17, n19, n20,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n190, n191, n192, n193, n194,
         n196, n197, n198, n200, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ps;

  DFFX1 \reg_b_reg[0]  ( .D(N66), .CLK(clk), .Q(reg_b[0]), .QN(n204) );
  DFFX1 \reg_b_reg[20]  ( .D(N86), .CLK(clk), .Q(reg_b[20]), .QN(n211) );
  DFFX1 \reg_a_reg[4]  ( .D(N30), .CLK(clk), .Q(result[4]), .QN(n203) );
  DFFX1 \reg_a_reg[1]  ( .D(N27), .CLK(clk), .Q(result[1]), .QN(n202) );
  DFFX1 \reg_a_reg[3]  ( .D(N29), .CLK(clk), .QN(n120) );
  DFFX2 \reg_a_reg[0]  ( .D(N26), .CLK(clk), .QN(n221) );
  DFFX1 \reg_a_reg[29]  ( .D(N55), .CLK(clk), .Q(result[29]), .QN(n156) );
  DFFX1 \reg_b_reg[9]  ( .D(N75), .CLK(clk), .Q(reg_b[9]), .QN(n157) );
  DFFX1 \reg_b_reg[25]  ( .D(N91), .CLK(clk), .Q(reg_b[25]), .QN(n174) );
  DFFX1 \reg_b_reg[21]  ( .D(N87), .CLK(clk), .Q(reg_b[21]), .QN(n172) );
  DFFX1 \reg_b_reg[14]  ( .D(N80), .CLK(clk), .Q(reg_b[14]), .QN(n171) );
  DFFX1 \reg_b_reg[17]  ( .D(N83), .CLK(clk), .Q(reg_b[17]), .QN(n166) );
  DFFX1 \reg_b_reg[13]  ( .D(N79), .CLK(clk), .Q(reg_b[13]), .QN(n165) );
  DFFX1 \reg_b_reg[19]  ( .D(N85), .CLK(clk), .Q(reg_b[19]), .QN(n178) );
  DFFX1 \reg_b_reg[15]  ( .D(N81), .CLK(clk), .Q(reg_b[15]), .QN(n168) );
  DFFX1 \reg_b_reg[11]  ( .D(N77), .CLK(clk), .Q(reg_b[11]), .QN(n167) );
  DFFX1 \reg_b_reg[27]  ( .D(N93), .CLK(clk), .Q(reg_b[27]), .QN(n175) );
  DFFX1 \reg_b_reg[23]  ( .D(N89), .CLK(clk), .Q(reg_b[23]), .QN(n173) );
  DFFX1 \reg_a_reg[30]  ( .D(N56), .CLK(clk), .Q(result[30]), .QN(n162) );
  DFFX1 \reg_a_reg[16]  ( .D(N42), .CLK(clk), .Q(result[16]), .QN(n140) );
  DFFX1 \reg_b_reg[26]  ( .D(N92), .CLK(clk), .Q(reg_b[26]), .QN(n177) );
  DFFX1 \reg_b_reg[22]  ( .D(N88), .CLK(clk), .Q(reg_b[22]), .QN(n164) );
  DFFX1 \reg_b_reg[28]  ( .D(N94), .CLK(clk), .Q(reg_b[28]), .QN(n155) );
  DFFX1 \reg_b_reg[24]  ( .D(N90), .CLK(clk), .Q(reg_b[24]), .QN(n163) );
  DFFX1 \reg_a_reg[13]  ( .D(N39), .CLK(clk), .Q(result[13]), .QN(n169) );
  DFFX1 \reg_a_reg[14]  ( .D(N40), .CLK(clk), .Q(result[14]), .QN(n134) );
  DFFX1 \reg_a_reg[18]  ( .D(N44), .CLK(clk), .Q(result[18]), .QN(n136) );
  DFFX1 \reg_a_reg[27]  ( .D(N53), .CLK(clk), .Q(result[27]), .QN(n158) );
  DFFX1 \reg_a_reg[25]  ( .D(N51), .CLK(clk), .Q(result[25]), .QN(n161) );
  DFFX1 \reg_a_reg[23]  ( .D(N49), .CLK(clk), .Q(result[23]), .QN(n159) );
  DFFX1 \reg_a_reg[21]  ( .D(N47), .CLK(clk), .Q(result[21]), .QN(n160) );
  DFFX1 \reg_a_reg[11]  ( .D(N37), .CLK(clk), .Q(result[11]), .QN(n180) );
  DFFX1 \reg_a_reg[17]  ( .D(N43), .CLK(clk), .Q(result[17]), .QN(n170) );
  DFFX1 \reg_a_reg[22]  ( .D(N48), .CLK(clk), .Q(result[22]), .QN(n176) );
  DFFARX1 \gcd_ps_reg[1]  ( .D(n71), .CLK(clk), .RSTB(reset_n), .Q(gcd_ps[1])
         );
  DFFARX1 \gcd_ps_reg[0]  ( .D(n72), .CLK(clk), .RSTB(reset_n), .Q(gcd_ps[0]), 
        .QN(n264) );
  DFFSSRX1 \reg_b_reg[4]  ( .SETB(1'b1), .RSTB(1'b1), .D(N70), .CLK(clk), .Q(
        n198), .QN(n88) );
  DFFX1 \reg_b_reg[8]  ( .D(N74), .CLK(clk), .Q(n73), .QN(n187) );
  DFFX1 \reg_b_reg[16]  ( .D(N82), .CLK(clk), .Q(reg_b[16]) );
  DFFX1 \reg_b_reg[7]  ( .D(N73), .CLK(clk), .Q(n77), .QN(n192) );
  DFFX1 \reg_b_reg[5]  ( .D(N71), .CLK(clk), .Q(n74), .QN(n190) );
  DFFX1 \reg_b_reg[10]  ( .D(N76), .CLK(clk), .Q(reg_b[10]) );
  DFFX1 \reg_b_reg[6]  ( .D(N72), .CLK(clk), .Q(reg_b[6]) );
  DFFX1 \reg_b_reg[29]  ( .D(N95), .CLK(clk), .Q(reg_b[29]) );
  DFFX1 \reg_b_reg[12]  ( .D(N78), .CLK(clk), .Q(reg_b[12]) );
  DFFX1 \reg_b_reg[2]  ( .D(N68), .CLK(clk), .Q(reg_b[2]), .QN(n329) );
  DFFX1 \reg_b_reg[31]  ( .D(N97), .CLK(clk), .Q(reg_b[31]) );
  DFFX1 \reg_b_reg[30]  ( .D(N96), .CLK(clk), .Q(reg_b[30]) );
  DFFX1 \reg_a_reg[7]  ( .D(N33), .CLK(clk), .QN(n188) );
  DFFX1 \reg_a_reg[9]  ( .D(N35), .CLK(clk), .QN(n194) );
  DFFX1 \reg_a_reg[6]  ( .D(N32), .CLK(clk), .Q(result[6]), .QN(n284) );
  DFFX1 \reg_a_reg[2]  ( .D(N28), .CLK(clk), .Q(result[2]), .QN(n196) );
  DFFX1 \reg_a_reg[28]  ( .D(N54), .CLK(clk), .Q(result[28]) );
  DFFX1 \reg_a_reg[26]  ( .D(N52), .CLK(clk), .Q(result[26]) );
  DFFX1 \reg_a_reg[24]  ( .D(N50), .CLK(clk), .Q(result[24]) );
  DFFX1 \reg_a_reg[20]  ( .D(N46), .CLK(clk), .Q(result[20]) );
  DFFX1 \reg_a_reg[19]  ( .D(N45), .CLK(clk), .Q(result[19]) );
  DFFX1 \reg_a_reg[12]  ( .D(N38), .CLK(clk), .Q(result[12]), .QN(n274) );
  DFFX1 \reg_a_reg[10]  ( .D(N36), .CLK(clk), .Q(result[10]), .QN(n271) );
  DFFX1 \reg_a_reg[8]  ( .D(N34), .CLK(clk), .Q(result[8]), .QN(n197) );
  DFFX1 \reg_a_reg[5]  ( .D(N31), .CLK(clk), .QN(n200) );
  DFFX1 \reg_a_reg[31]  ( .D(N57), .CLK(clk), .Q(result[31]), .QN(n318) );
  DFFX1 \reg_b_reg[18]  ( .D(N84), .CLK(clk), .Q(reg_b[18]), .QN(n269) );
  DFFX1 \reg_b_reg[3]  ( .D(N69), .CLK(clk), .Q(n89), .QN(n191) );
  DFFX1 \reg_b_reg[1]  ( .D(N67), .CLK(clk), .QN(n119) );
  DFFX2 \reg_a_reg[15]  ( .D(N41), .CLK(clk), .Q(result[15]) );
  NAND2X1 U135 ( .IN1(n87), .IN2(n347), .QN(n98) );
  XOR3X2 U136 ( .IN1(result[11]), .IN2(reg_b[11]), .IN3(n85), .Q(n379) );
  NAND2X4 U137 ( .IN1(n167), .IN2(result[11]), .QN(n380) );
  XOR3X2 U138 ( .IN1(result[15]), .IN2(reg_b[15]), .IN3(n133), .Q(n398) );
  NAND2X4 U139 ( .IN1(n168), .IN2(result[15]), .QN(n399) );
  NAND2X2 U140 ( .IN1(n287), .IN2(n288), .QN(n392) );
  NOR2X1 U141 ( .IN1(n372), .IN2(n280), .QN(n286) );
  NOR2X0 U142 ( .IN1(reg_b[2]), .IN2(n196), .QN(n181) );
  OAI21X1 U143 ( .IN1(result[2]), .IN2(n329), .IN3(n324), .QN(n109) );
  NAND2X2 U144 ( .IN1(n121), .IN2(n84), .QN(n373) );
  NAND2X2 U145 ( .IN1(n285), .IN2(n345), .QN(n121) );
  INVX2 U146 ( .IN(n402), .QN(n291) );
  NAND2X0 U147 ( .IN1(n297), .IN2(n296), .QN(n298) );
  NOR2X0 U148 ( .IN1(n293), .IN2(n292), .QN(n297) );
  NAND2X0 U149 ( .IN1(n411), .IN2(n295), .QN(n296) );
  INVX0 U150 ( .IN(n419), .QN(n293) );
  INVX0 U151 ( .IN(n387), .QN(n270) );
  INVX0 U152 ( .IN(n357), .QN(n278) );
  NAND2X2 U153 ( .IN1(n190), .IN2(result[5]), .QN(n351) );
  NOR2X0 U154 ( .IN1(reg_b[16]), .IN2(n140), .QN(n186) );
  AND2X1 U155 ( .IN1(n154), .IN2(n109), .Q(n348) );
  NAND2X2 U156 ( .IN1(n262), .IN2(result[9]), .QN(n228) );
  NAND2X0 U157 ( .IN1(n215), .IN2(reg_b[9]), .QN(n106) );
  NAND2X0 U158 ( .IN1(n166), .IN2(result[17]), .QN(n407) );
  INVX2 U159 ( .IN(n194), .QN(result[9]) );
  OAI21X1 U160 ( .IN1(result[2]), .IN2(n329), .IN3(n324), .QN(n345) );
  NAND2X0 U161 ( .IN1(n380), .IN2(n375), .QN(n280) );
  INVX0 U162 ( .IN(n279), .QN(n272) );
  NAND2X0 U163 ( .IN1(n399), .IN2(n394), .QN(n289) );
  AO221X1 U164 ( .IN1(n290), .IN2(n395), .IN3(reg_b[16]), .IN4(n140), .IN5(
        n182), .Q(n402) );
  INVX0 U165 ( .IN(start), .QN(n321) );
  OAI21X1 U166 ( .IN1(result[18]), .IN2(n269), .IN3(n406), .QN(n415) );
  NOR2X2 U167 ( .IN1(n112), .IN2(n114), .QN(n229) );
  INVX0 U168 ( .IN(n102), .QN(n384) );
  OA21X1 U169 ( .IN1(n16), .IN2(n143), .IN3(n323), .Q(n206) );
  OR2X1 U170 ( .IN1(result[3]), .IN2(n191), .Q(n340) );
  INVX0 U171 ( .IN(n323), .QN(n485) );
  INVX0 U172 ( .IN(n322), .QN(n487) );
  AND2X1 U173 ( .IN1(n478), .IN2(n477), .Q(n479) );
  INVX0 U174 ( .IN(n108), .QN(n354) );
  NAND2X0 U175 ( .IN1(n157), .IN2(result[9]), .QN(n368) );
  AND2X1 U176 ( .IN1(n363), .IN2(n108), .Q(n366) );
  XOR3X1 U177 ( .IN1(reg_b[6]), .IN2(result[6]), .IN3(n352), .Q(n353) );
  INVX0 U178 ( .IN(a_in[7]), .QN(n104) );
  AND2X1 U179 ( .IN1(n374), .IN2(n108), .Q(n377) );
  NAND2X0 U180 ( .IN1(n165), .IN2(result[13]), .QN(n387) );
  AND2X1 U181 ( .IN1(n393), .IN2(n102), .Q(n396) );
  INVX2 U182 ( .IN(n223), .QN(n224) );
  OAI21X1 U183 ( .IN1(n469), .IN2(n213), .IN3(n468), .QN(n478) );
  AND2X1 U184 ( .IN1(n462), .IN2(n463), .Q(n213) );
  NAND2X2 U185 ( .IN1(n486), .IN2(n206), .QN(n474) );
  INVX0 U186 ( .IN(n97), .QN(n488) );
  INVX2 U187 ( .IN(n119), .QN(n193) );
  OR2X1 U188 ( .IN1(n89), .IN2(n281), .Q(n341) );
  NBUFFX2 U189 ( .IN(n490), .Q(n263) );
  INVX0 U190 ( .IN(n109), .QN(n336) );
  INVX4 U191 ( .IN(n120), .QN(result[3]) );
  INVX2 U192 ( .IN(n200), .QN(result[5]) );
  NAND2X0 U193 ( .IN1(n232), .IN2(n233), .QN(n437) );
  NOR2X0 U194 ( .IN1(n327), .IN2(n326), .QN(n335) );
  NOR2X0 U195 ( .IN1(n333), .IN2(n332), .QN(n334) );
  NAND2X1 U196 ( .IN1(n81), .IN2(n94), .QN(N35) );
  XOR3X1 U197 ( .IN1(result[25]), .IN2(reg_b[25]), .IN3(n128), .Q(n444) );
  XOR3X1 U198 ( .IN1(result[27]), .IN2(reg_b[27]), .IN3(n148), .Q(n454) );
  XOR3X1 U199 ( .IN1(reg_b[18]), .IN2(n136), .IN3(n137), .Q(n410) );
  NAND2X0 U200 ( .IN1(n261), .IN2(result[13]), .QN(n218) );
  INVX1 U201 ( .IN(n225), .QN(n209) );
  INVX1 U202 ( .IN(n330), .QN(n205) );
  NOR2X0 U203 ( .IN1(result[19]), .IN2(n178), .QN(n78) );
  AND2X1 U204 ( .IN1(n160), .IN2(reg_b[21]), .Q(n79) );
  OR3X1 U205 ( .IN1(n321), .IN2(gcd_ps[0]), .IN3(gcd_ps[1]), .Q(n322) );
  NOR2X0 U206 ( .IN1(reg_b[31]), .IN2(n318), .QN(n80) );
  AND2X1 U207 ( .IN1(n105), .IN2(n106), .Q(n81) );
  AOI22X1 U208 ( .IN1(a_in[6]), .IN2(n225), .IN3(n215), .IN4(reg_b[6]), .QN(
        n82) );
  AOI22X1 U209 ( .IN1(a_in[13]), .IN2(n225), .IN3(n215), .IN4(reg_b[13]), .QN(
        n83) );
  AND3X1 U210 ( .IN1(n98), .IN2(n99), .IN3(n100), .Q(n84) );
  OA21X1 U211 ( .IN1(n377), .IN2(n376), .IN3(n375), .Q(n85) );
  OA21X1 U212 ( .IN1(n366), .IN2(n365), .IN3(n364), .Q(n86) );
  AND2X1 U213 ( .IN1(n351), .IN2(n346), .Q(n87) );
  INVX2 U214 ( .IN(n188), .QN(result[7]) );
  NOR2X0 U215 ( .IN1(n415), .IN2(n299), .QN(n90) );
  AOI22X1 U216 ( .IN1(a_in[0]), .IN2(n225), .IN3(n489), .IN4(reg_b[0]), .QN(
        n91) );
  AND2X1 U217 ( .IN1(n110), .IN2(n111), .Q(n92) );
  AND2X1 U218 ( .IN1(n217), .IN2(n218), .Q(n93) );
  AND2X1 U219 ( .IN1(n227), .IN2(n228), .Q(n94) );
  AND2X1 U220 ( .IN1(n123), .IN2(n124), .Q(n95) );
  INVX4 U221 ( .IN(n474), .QN(n490) );
  NBUFFX2 U222 ( .IN(n490), .Q(n257) );
  INVX0 U223 ( .IN(n215), .QN(n216) );
  INVX8 U224 ( .IN(n337), .QN(n215) );
  INVX2 U225 ( .IN(n223), .QN(n225) );
  NOR2X4 U227 ( .IN1(result[0]), .IN2(n204), .QN(n97) );
  NAND2X0 U228 ( .IN1(reg_b[6]), .IN2(n284), .QN(n99) );
  INVX0 U229 ( .IN(n153), .QN(n100) );
  OAI21X1 U230 ( .IN1(result[4]), .IN2(n88), .IN3(n340), .QN(n347) );
  INVX4 U231 ( .IN(n101), .QN(n472) );
  NOR2X2 U232 ( .IN1(n206), .IN2(n328), .QN(n101) );
  MUX21X1 U233 ( .IN1(n470), .IN2(n471), .S(n478), .Q(n473) );
  INVX4 U234 ( .IN(n328), .QN(n486) );
  NAND2X0 U235 ( .IN1(n287), .IN2(n288), .QN(n102) );
  NAND2X0 U236 ( .IN1(n178), .IN2(result[19]), .QN(n419) );
  OA22X1 U237 ( .IN1(n104), .IN2(n209), .IN3(n337), .IN4(n192), .Q(n103) );
  NAND2X2 U238 ( .IN1(n83), .IN2(n93), .QN(N39) );
  NAND2X1 U239 ( .IN1(n492), .IN2(n385), .QN(n217) );
  NAND2X0 U240 ( .IN1(a_in[9]), .IN2(n225), .QN(n105) );
  NAND2X1 U241 ( .IN1(n492), .IN2(n367), .QN(n227) );
  NAND2X2 U242 ( .IN1(n82), .IN2(n92), .QN(N32) );
  NAND2X1 U243 ( .IN1(n492), .IN2(n353), .QN(n110) );
  OR2X1 U244 ( .IN1(n16), .IN2(n143), .Q(n107) );
  NAND2X1 U245 ( .IN1(n107), .IN2(n323), .QN(n330) );
  DELLN1X2 U246 ( .IN(n373), .Q(n108) );
  NAND2X0 U247 ( .IN1(n263), .IN2(result[6]), .QN(n111) );
  AND3X1 U248 ( .IN1(n392), .IN2(n290), .IN3(n393), .Q(n112) );
  OR2X1 U249 ( .IN1(n270), .IN2(n183), .Q(n391) );
  NOR3X0 U250 ( .IN1(n391), .IN2(n289), .IN3(n384), .QN(n113) );
  OA21X1 U251 ( .IN1(n457), .IN2(n148), .IN3(n456), .Q(n458) );
  NAND2X1 U252 ( .IN1(n291), .IN2(n90), .QN(n114) );
  NAND2X0 U253 ( .IN1(n492), .IN2(n491), .QN(n115) );
  NAND2X0 U254 ( .IN1(n257), .IN2(result[0]), .QN(n116) );
  NAND3X0 U255 ( .IN1(n115), .IN2(n116), .IN3(n91), .QN(N26) );
  NAND2X2 U256 ( .IN1(n215), .IN2(reg_b[24]), .QN(n233) );
  INVX1 U257 ( .IN(n117), .QN(n226) );
  NAND2X4 U258 ( .IN1(n122), .IN2(n95), .QN(n376) );
  NAND2X4 U259 ( .IN1(n272), .IN2(n365), .QN(n122) );
  INVX0 U260 ( .IN(n185), .QN(n124) );
  NAND2X4 U261 ( .IN1(n273), .IN2(n376), .QN(n276) );
  NOR2X4 U262 ( .IN1(n302), .IN2(n125), .QN(n126) );
  INVX8 U263 ( .IN(n223), .QN(n117) );
  INVX8 U264 ( .IN(n223), .QN(n118) );
  NOR2X4 U265 ( .IN1(n146), .IN2(n300), .QN(n302) );
  INVX0 U266 ( .IN(n126), .QN(n150) );
  NAND2X2 U267 ( .IN1(n276), .IN2(n275), .QN(n277) );
  OAI21X1 U268 ( .IN1(result[8]), .IN2(n187), .IN3(n356), .QN(n365) );
  NAND2X0 U269 ( .IN1(n170), .IN2(reg_b[17]), .QN(n406) );
  NAND2X2 U270 ( .IN1(n169), .IN2(reg_b[13]), .QN(n386) );
  NAND2X0 U271 ( .IN1(reg_b[10]), .IN2(n271), .QN(n123) );
  OR2X1 U272 ( .IN1(n301), .IN2(n79), .Q(n125) );
  NOR2X0 U273 ( .IN1(n268), .IN2(n315), .QN(n317) );
  NAND2X0 U274 ( .IN1(n440), .IN2(n446), .QN(n307) );
  NAND2X0 U275 ( .IN1(n430), .IN2(n434), .QN(n303) );
  NBUFFX2 U276 ( .IN(n487), .Q(n249) );
  NOR2X1 U277 ( .IN1(reg_b[6]), .IN2(n284), .QN(n184) );
  NAND2X0 U278 ( .IN1(n173), .IN2(result[23]), .QN(n434) );
  NAND2X0 U279 ( .IN1(n211), .IN2(result[20]), .QN(n423) );
  NAND2X0 U280 ( .IN1(n172), .IN2(result[21]), .QN(n427) );
  NAND2X1 U281 ( .IN1(n171), .IN2(result[14]), .QN(n394) );
  INVX2 U282 ( .IN(n289), .QN(n290) );
  NAND2X0 U283 ( .IN1(n269), .IN2(result[18]), .QN(n414) );
  AND2X1 U284 ( .IN1(n176), .IN2(reg_b[22]), .Q(n301) );
  NAND2X2 U285 ( .IN1(n368), .IN2(n364), .QN(n279) );
  INVX0 U286 ( .IN(n280), .QN(n273) );
  NOR2X0 U287 ( .IN1(n186), .IN2(n403), .QN(n127) );
  NOR2X0 U288 ( .IN1(n442), .IN2(n441), .QN(n128) );
  NOR2X0 U289 ( .IN1(n146), .IN2(n424), .QN(n129) );
  NOR2X0 U290 ( .IN1(n354), .IN2(n184), .QN(n130) );
  NOR2X0 U291 ( .IN1(n336), .IN2(n181), .QN(n131) );
  OA21X1 U292 ( .IN1(n416), .IN2(n415), .IN3(n414), .Q(n132) );
  OA21X1 U293 ( .IN1(n396), .IN2(n395), .IN3(n394), .Q(n133) );
  INVX0 U294 ( .IN(result[3]), .QN(n281) );
  NOR2X0 U295 ( .IN1(result[24]), .IN2(n163), .QN(n304) );
  NOR2X0 U296 ( .IN1(result[26]), .IN2(n177), .QN(n308) );
  NOR2X0 U297 ( .IN1(result[28]), .IN2(n155), .QN(n312) );
  NOR2X0 U298 ( .IN1(result[15]), .IN2(n168), .QN(n182) );
  NOR2X0 U299 ( .IN1(result[20]), .IN2(n211), .QN(n299) );
  XOR3X1 U300 ( .IN1(n134), .IN2(reg_b[14]), .IN3(n135), .Q(n390) );
  OAI21X1 U301 ( .IN1(n388), .IN2(n152), .IN3(n387), .QN(n135) );
  OAI21X1 U302 ( .IN1(n408), .IN2(n127), .IN3(n407), .QN(n137) );
  XOR3X1 U303 ( .IN1(n164), .IN2(result[22]), .IN3(n138), .Q(n429) );
  OAI21X1 U304 ( .IN1(n79), .IN2(n129), .IN3(n427), .QN(n138) );
  XOR3X1 U305 ( .IN1(n177), .IN2(result[26]), .IN3(n139), .Q(n449) );
  OAI21X1 U306 ( .IN1(n447), .IN2(n128), .IN3(n446), .QN(n139) );
  XOR3X1 U307 ( .IN1(n140), .IN2(reg_b[16]), .IN3(n141), .Q(n401) );
  OAI21X1 U308 ( .IN1(n182), .IN2(n133), .IN3(n399), .QN(n141) );
  OA21X2 U309 ( .IN1(n480), .IN2(n479), .IN3(n80), .Q(n482) );
  XOR3X1 U310 ( .IN1(n203), .IN2(n198), .IN3(n142), .Q(n344) );
  OAI21X1 U311 ( .IN1(n342), .IN2(n131), .IN3(n341), .QN(n142) );
  OR2X1 U312 ( .IN1(reg_b[10]), .IN2(n271), .Q(n375) );
  NOR2X4 U313 ( .IN1(n277), .IN2(n179), .QN(n288) );
  NBUFFX2 U314 ( .IN(n485), .Q(n240) );
  NBUFFX2 U315 ( .IN(n490), .Q(n259) );
  NBUFFX2 U316 ( .IN(n490), .Q(n261) );
  NBUFFX2 U317 ( .IN(n490), .Q(n262) );
  NBUFFX2 U318 ( .IN(n490), .Q(n258) );
  NAND2X4 U319 ( .IN1(n323), .IN2(n322), .QN(n328) );
  OR2X1 U320 ( .IN1(n362), .IN2(n279), .Q(n372) );
  INVX0 U321 ( .IN(n356), .QN(n358) );
  INVX0 U322 ( .IN(n340), .QN(n342) );
  OR2X1 U323 ( .IN1(n77), .IN2(n188), .Q(n357) );
  NOR2X0 U324 ( .IN1(n16), .IN2(n80), .QN(n319) );
  OR2X1 U325 ( .IN1(n294), .IN2(n186), .Q(n411) );
  INVX0 U326 ( .IN(n407), .QN(n294) );
  OR2X1 U327 ( .IN1(n278), .IN2(n184), .Q(n362) );
  OR2X1 U328 ( .IN1(n113), .IN2(n402), .Q(n412) );
  NOR2X0 U329 ( .IN1(n266), .IN2(n265), .QN(n268) );
  XOR3X1 U330 ( .IN1(result[7]), .IN2(n77), .IN3(n130), .Q(n355) );
  INVX0 U331 ( .IN(n391), .QN(n393) );
  AND2X1 U332 ( .IN1(n144), .IN2(n145), .Q(n143) );
  NOR4X0 U333 ( .IN1(n64), .IN2(n63), .IN3(n66), .IN4(n65), .QN(n144) );
  NOR4X0 U334 ( .IN1(n68), .IN2(n67), .IN3(n70), .IN4(n69), .QN(n145) );
  OR2X1 U335 ( .IN1(n73), .IN2(n197), .Q(n364) );
  AND2X1 U336 ( .IN1(result[2]), .IN2(n260), .Q(n327) );
  NAND2X0 U337 ( .IN1(n423), .IN2(n427), .QN(n300) );
  NOR2X4 U338 ( .IN1(n147), .IN2(n78), .QN(n146) );
  NOR2X4 U339 ( .IN1(n229), .IN2(n230), .QN(n147) );
  OR2X1 U340 ( .IN1(result[7]), .IN2(n192), .Q(n356) );
  NAND2X0 U341 ( .IN1(n476), .IN2(n468), .QN(n265) );
  NAND2X0 U342 ( .IN1(n451), .IN2(n456), .QN(n311) );
  INVX0 U343 ( .IN(n463), .QN(n266) );
  AND2X1 U344 ( .IN1(n450), .IN2(n451), .Q(n148) );
  AND2X1 U345 ( .IN1(n150), .IN2(n430), .Q(n149) );
  NBUFFX2 U346 ( .IN(n487), .Q(n252) );
  NBUFFX2 U347 ( .IN(n487), .Q(n253) );
  NBUFFX2 U348 ( .IN(n487), .Q(n254) );
  NBUFFX2 U349 ( .IN(n487), .Q(n255) );
  NBUFFX2 U350 ( .IN(n487), .Q(n251) );
  NBUFFX2 U351 ( .IN(n487), .Q(n256) );
  NBUFFX2 U352 ( .IN(n487), .Q(n250) );
  NAND2X1 U353 ( .IN1(n335), .IN2(n334), .QN(N28) );
  AND2X1 U354 ( .IN1(n461), .IN2(n468), .Q(n465) );
  INVX0 U355 ( .IN(n15), .QN(n494) );
  INVX0 U356 ( .IN(n461), .QN(n469) );
  INVX0 U357 ( .IN(n362), .QN(n363) );
  OA21X1 U358 ( .IN1(n348), .IN2(n347), .IN3(n346), .Q(n151) );
  INVX0 U359 ( .IN(n372), .QN(n374) );
  INVX0 U360 ( .IN(n20), .QN(done) );
  INVX0 U361 ( .IN(n415), .QN(n295) );
  AND2X1 U362 ( .IN1(n413), .IN2(n412), .Q(n416) );
  INVX0 U363 ( .IN(n411), .QN(n413) );
  INVX0 U364 ( .IN(n440), .QN(n441) );
  NOR2X0 U365 ( .IN1(n384), .IN2(n183), .QN(n152) );
  INVX0 U366 ( .IN(n423), .QN(n424) );
  INVX0 U367 ( .IN(n412), .QN(n403) );
  NOR2X0 U368 ( .IN1(result[5]), .IN2(n190), .QN(n153) );
  INVX0 U369 ( .IN(n414), .QN(n292) );
  NOR2X4 U370 ( .IN1(n282), .IN2(n181), .QN(n154) );
  AND2X1 U371 ( .IN1(n477), .IN2(n476), .Q(n471) );
  INVX0 U372 ( .IN(n433), .QN(n435) );
  INVX0 U373 ( .IN(n445), .QN(n447) );
  INVX0 U374 ( .IN(n455), .QN(n457) );
  INVX0 U375 ( .IN(n406), .QN(n408) );
  INVX0 U376 ( .IN(n386), .QN(n388) );
  NAND2X0 U377 ( .IN1(n155), .IN2(result[28]), .QN(n463) );
  INVX0 U378 ( .IN(a_in[2]), .QN(n331) );
  AO221X1 U379 ( .IN1(start), .IN2(n264), .IN3(n143), .IN4(n493), .IN5(n19), 
        .Q(n15) );
  INVX0 U380 ( .IN(n16), .QN(n493) );
  NAND2X0 U381 ( .IN1(reset_n), .IN2(n20), .QN(n19) );
  NAND2X0 U382 ( .IN1(n156), .IN2(reg_b[29]), .QN(n461) );
  NAND2X0 U383 ( .IN1(gcd_ps[1]), .IN2(n264), .QN(n20) );
  AO221X1 U384 ( .IN1(n469), .IN2(n476), .IN3(reg_b[31]), .IN4(n318), .IN5(
        n267), .Q(n315) );
  INVX0 U385 ( .IN(n477), .QN(n267) );
  OR2X1 U386 ( .IN1(reg_b[30]), .IN2(n162), .Q(n476) );
  AO222X1 U387 ( .IN1(b_in[31]), .IN2(n256), .IN3(n248), .IN4(reg_b[31]), 
        .IN5(n236), .IN6(result[31]), .Q(N97) );
  AO222X1 U388 ( .IN1(b_in[16]), .IN2(n252), .IN3(n242), .IN4(reg_b[16]), 
        .IN5(n236), .IN6(result[16]), .Q(N82) );
  AO222X1 U389 ( .IN1(b_in[6]), .IN2(n250), .IN3(n244), .IN4(reg_b[6]), .IN5(
        n240), .IN6(result[6]), .Q(N72) );
  AO222X1 U390 ( .IN1(b_in[10]), .IN2(n251), .IN3(n243), .IN4(reg_b[10]), 
        .IN5(n238), .IN6(result[10]), .Q(N76) );
  AO222X1 U391 ( .IN1(b_in[12]), .IN2(n251), .IN3(n246), .IN4(reg_b[12]), 
        .IN5(n239), .IN6(result[12]), .Q(N78) );
  AO222X1 U392 ( .IN1(b_in[21]), .IN2(n254), .IN3(n248), .IN4(reg_b[21]), 
        .IN5(n240), .IN6(result[21]), .Q(N87) );
  AO222X1 U393 ( .IN1(b_in[27]), .IN2(n255), .IN3(n248), .IN4(reg_b[27]), 
        .IN5(n237), .IN6(result[27]), .Q(N93) );
  AO222X1 U394 ( .IN1(b_in[11]), .IN2(n251), .IN3(n247), .IN4(reg_b[11]), 
        .IN5(n237), .IN6(result[11]), .Q(N77) );
  AO222X1 U395 ( .IN1(b_in[13]), .IN2(n252), .IN3(n245), .IN4(reg_b[13]), 
        .IN5(n236), .IN6(result[13]), .Q(N79) );
  AO222X1 U396 ( .IN1(b_in[23]), .IN2(n254), .IN3(n245), .IN4(reg_b[23]), 
        .IN5(n237), .IN6(result[23]), .Q(N89) );
  AO222X1 U397 ( .IN1(b_in[15]), .IN2(n252), .IN3(n243), .IN4(reg_b[15]), 
        .IN5(n238), .IN6(result[15]), .Q(N81) );
  AO222X1 U398 ( .IN1(b_in[17]), .IN2(n253), .IN3(n241), .IN4(reg_b[17]), 
        .IN5(n239), .IN6(result[17]), .Q(N83) );
  AO222X1 U399 ( .IN1(b_in[18]), .IN2(n253), .IN3(n242), .IN4(reg_b[18]), 
        .IN5(n240), .IN6(result[18]), .Q(N84) );
  AO222X1 U400 ( .IN1(b_in[19]), .IN2(n253), .IN3(n241), .IN4(reg_b[19]), 
        .IN5(n235), .IN6(result[19]), .Q(N85) );
  AO222X1 U401 ( .IN1(b_in[25]), .IN2(n255), .IN3(n243), .IN4(reg_b[25]), 
        .IN5(n238), .IN6(result[25]), .Q(N91) );
  AO222X1 U402 ( .IN1(b_in[14]), .IN2(n252), .IN3(n244), .IN4(reg_b[14]), 
        .IN5(n235), .IN6(result[14]), .Q(N80) );
  AO222X1 U403 ( .IN1(b_in[30]), .IN2(n256), .IN3(n241), .IN4(reg_b[30]), 
        .IN5(n234), .IN6(result[30]), .Q(N96) );
  AO222X1 U404 ( .IN1(b_in[26]), .IN2(n255), .IN3(n248), .IN4(reg_b[26]), 
        .IN5(n234), .IN6(result[26]), .Q(N92) );
  AO222X1 U405 ( .IN1(b_in[28]), .IN2(n255), .IN3(n248), .IN4(reg_b[28]), 
        .IN5(n240), .IN6(result[28]), .Q(N94) );
  AO222X1 U406 ( .IN1(b_in[22]), .IN2(n254), .IN3(n246), .IN4(reg_b[22]), 
        .IN5(n234), .IN6(result[22]), .Q(N88) );
  AO222X1 U407 ( .IN1(b_in[24]), .IN2(n254), .IN3(n244), .IN4(reg_b[24]), 
        .IN5(n235), .IN6(result[24]), .Q(N90) );
  AO222X1 U408 ( .IN1(b_in[20]), .IN2(n253), .IN3(n244), .IN4(reg_b[20]), 
        .IN5(n235), .IN6(result[20]), .Q(N86) );
  AO222X1 U409 ( .IN1(b_in[1]), .IN2(n256), .IN3(n247), .IN4(n193), .IN5(n239), 
        .IN6(result[1]), .Q(N67) );
  OR4X1 U410 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(
        reg_b[16]), .Q(n69) );
  OR4X1 U411 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n65) );
  OR4X1 U412 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n66) );
  OR4X1 U413 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n67) );
  OR4X1 U414 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(n193), 
        .Q(n68) );
  NAND2X0 U415 ( .IN1(n158), .IN2(reg_b[27]), .QN(n455) );
  NAND2X0 U416 ( .IN1(n159), .IN2(reg_b[23]), .QN(n433) );
  NAND2X0 U417 ( .IN1(n161), .IN2(reg_b[25]), .QN(n445) );
  NAND2X0 U418 ( .IN1(n162), .IN2(reg_b[30]), .QN(n477) );
  NAND2X0 U419 ( .IN1(n163), .IN2(result[24]), .QN(n440) );
  NAND2X0 U420 ( .IN1(n164), .IN2(result[22]), .QN(n430) );
  AO22X1 U421 ( .IN1(n494), .IN2(gcd_ps[1]), .IN3(n14), .IN4(n15), .Q(n71) );
  NAND2X0 U422 ( .IN1(n16), .IN2(reset_n), .QN(n14) );
  XOR3X1 U423 ( .IN1(n193), .IN2(result[1]), .IN3(n97), .Q(n484) );
  XOR3X1 U424 ( .IN1(result[21]), .IN2(reg_b[21]), .IN3(n129), .Q(n426) );
  INVX0 U425 ( .IN(n209), .QN(n208) );
  OR2X1 U426 ( .IN1(reg_b[29]), .IN2(n156), .Q(n468) );
  XOR3X1 U427 ( .IN1(result[17]), .IN2(reg_b[17]), .IN3(n127), .Q(n405) );
  XOR3X1 U428 ( .IN1(result[3]), .IN2(n89), .IN3(n131), .Q(n339) );
  XOR3X1 U429 ( .IN1(result[5]), .IN2(n74), .IN3(n151), .Q(n350) );
  XOR3X1 U430 ( .IN1(result[23]), .IN2(reg_b[23]), .IN3(n149), .Q(n432) );
  XOR3X1 U431 ( .IN1(result[10]), .IN2(reg_b[10]), .IN3(n369), .Q(n371) );
  OA21X1 U432 ( .IN1(n185), .IN2(n86), .IN3(n368), .Q(n369) );
  INVX0 U433 ( .IN(n476), .QN(n480) );
  XOR3X1 U434 ( .IN1(result[8]), .IN2(n73), .IN3(n359), .Q(n361) );
  OA21X1 U435 ( .IN1(n358), .IN2(n130), .IN3(n357), .Q(n359) );
  XOR3X1 U436 ( .IN1(result[19]), .IN2(reg_b[19]), .IN3(n132), .Q(n418) );
  OA21X1 U437 ( .IN1(n153), .IN2(n151), .IN3(n351), .Q(n352) );
  XOR3X1 U438 ( .IN1(reg_b[12]), .IN2(result[12]), .IN3(n381), .Q(n383) );
  OA21X1 U439 ( .IN1(n179), .IN2(n85), .IN3(n380), .Q(n381) );
  INVX0 U440 ( .IN(a_in[20]), .QN(n210) );
  XOR3X1 U441 ( .IN1(result[2]), .IN2(n324), .IN3(reg_b[2]), .Q(n325) );
  XOR3X1 U442 ( .IN1(result[9]), .IN2(reg_b[9]), .IN3(n86), .Q(n367) );
  XOR3X1 U443 ( .IN1(result[13]), .IN2(reg_b[13]), .IN3(n152), .Q(n385) );
  NAND2X0 U444 ( .IN1(n174), .IN2(result[25]), .QN(n446) );
  NAND2X0 U445 ( .IN1(n175), .IN2(result[27]), .QN(n456) );
  XOR3X1 U446 ( .IN1(reg_b[20]), .IN2(result[20]), .IN3(n420), .Q(n422) );
  OA21X1 U447 ( .IN1(n78), .IN2(n132), .IN3(n419), .Q(n420) );
  INVX0 U448 ( .IN(n226), .QN(n212) );
  MUX21X1 U449 ( .IN1(n465), .IN2(n464), .S(n213), .Q(n466) );
  XOR3X1 U450 ( .IN1(reg_b[24]), .IN2(result[24]), .IN3(n436), .Q(n438) );
  OA21X1 U451 ( .IN1(n435), .IN2(n149), .IN3(n434), .Q(n436) );
  INVX4 U452 ( .IN(n221), .QN(result[0]) );
  NAND2X0 U453 ( .IN1(reg_b[12]), .IN2(n274), .QN(n275) );
  OAI21X1 U454 ( .IN1(result[14]), .IN2(n171), .IN3(n386), .QN(n395) );
  OAI22X1 U455 ( .IN1(n264), .IN2(n15), .IN3(n494), .IN4(n17), .QN(n72) );
  OA21X1 U456 ( .IN1(gcd_ps[1]), .IN2(gcd_ps[0]), .IN3(reset_n), .Q(n17) );
  NAND2X0 U457 ( .IN1(n177), .IN2(result[26]), .QN(n451) );
  OR2X1 U458 ( .IN1(n264), .IN2(gcd_ps[1]), .Q(n16) );
  AND2X1 U459 ( .IN1(n180), .IN2(reg_b[11]), .Q(n179) );
  NOR2X0 U460 ( .IN1(reg_b[12]), .IN2(n274), .QN(n183) );
  NOR2X0 U461 ( .IN1(result[9]), .IN2(n157), .QN(n185) );
  XOR2X1 U462 ( .IN1(result[30]), .IN2(reg_b[30]), .Q(n470) );
  AO222X1 U463 ( .IN1(b_in[29]), .IN2(n256), .IN3(n247), .IN4(reg_b[29]), 
        .IN5(n234), .IN6(result[29]), .Q(N95) );
  XOR2X1 U464 ( .IN1(result[29]), .IN2(reg_b[29]), .Q(n464) );
  INVX4 U465 ( .IN(n439), .QN(n442) );
  AND2X1 U466 ( .IN1(n193), .IN2(n202), .Q(n283) );
  AO222X1 U467 ( .IN1(b_in[2]), .IN2(n249), .IN3(n247), .IN4(reg_b[2]), .IN5(
        n240), .IN6(result[2]), .Q(N68) );
  AO222X1 U468 ( .IN1(b_in[9]), .IN2(n251), .IN3(n241), .IN4(reg_b[9]), .IN5(
        n240), .IN6(result[9]), .Q(N75) );
  AO222X1 U469 ( .IN1(b_in[8]), .IN2(n250), .IN3(n242), .IN4(n73), .IN5(n240), 
        .IN6(result[8]), .Q(N74) );
  OR4X1 U470 ( .IN1(reg_b[6]), .IN2(n77), .IN3(n73), .IN4(reg_b[9]), .Q(n63)
         );
  AO222X1 U471 ( .IN1(b_in[7]), .IN2(n250), .IN3(n243), .IN4(n77), .IN5(n240), 
        .IN6(result[7]), .Q(N73) );
  OR2X2 U472 ( .IN1(n198), .IN2(n203), .Q(n346) );
  XOR3X1 U473 ( .IN1(reg_b[28]), .IN2(result[28]), .IN3(n458), .Q(n460) );
  OAI21X1 U474 ( .IN1(reg_b[0]), .IN2(n221), .IN3(n488), .QN(n491) );
  AO222X1 U475 ( .IN1(b_in[5]), .IN2(n250), .IN3(n245), .IN4(n74), .IN5(n236), 
        .IN6(result[5]), .Q(N71) );
  OR4X1 U476 ( .IN1(reg_b[31]), .IN2(n89), .IN3(n198), .IN4(n74), .Q(n64) );
  AO222X1 U477 ( .IN1(b_in[3]), .IN2(n249), .IN3(n246), .IN4(n89), .IN5(n238), 
        .IN6(result[3]), .Q(N69) );
  AND2X1 U478 ( .IN1(n87), .IN2(n154), .Q(n285) );
  INVX8 U479 ( .IN(n207), .QN(n337) );
  INVX4 U480 ( .IN(n450), .QN(n452) );
  NOR2X4 U481 ( .IN1(n486), .IN2(n205), .QN(n207) );
  INVX16 U482 ( .IN(n337), .QN(n489) );
  NBUFFX2 U483 ( .IN(n485), .Q(n239) );
  NBUFFX2 U484 ( .IN(n485), .Q(n238) );
  NBUFFX2 U485 ( .IN(n485), .Q(n237) );
  NBUFFX2 U486 ( .IN(n485), .Q(n236) );
  NBUFFX2 U487 ( .IN(n485), .Q(n235) );
  NBUFFX2 U488 ( .IN(n485), .Q(n234) );
  OAI22X1 U489 ( .IN1(n210), .IN2(n223), .IN3(n337), .IN4(n211), .QN(n421) );
  NBUFFX2 U490 ( .IN(n490), .Q(n260) );
  INVX8 U491 ( .IN(n214), .QN(n223) );
  INVX16 U492 ( .IN(n472), .QN(n492) );
  NOR2X4 U493 ( .IN1(n486), .IN2(n330), .QN(n214) );
  NAND2X0 U494 ( .IN1(n492), .IN2(n355), .QN(n219) );
  NAND2X0 U495 ( .IN1(n263), .IN2(result[7]), .QN(n220) );
  NAND3X0 U496 ( .IN1(n219), .IN2(n220), .IN3(n103), .QN(N33) );
  NOR2X0 U497 ( .IN1(n325), .IN2(n472), .QN(n326) );
  OAI22X1 U498 ( .IN1(n156), .IN2(n474), .IN3(n466), .IN4(n472), .QN(n467) );
  OAI22X1 U499 ( .IN1(n162), .IN2(n474), .IN3(n473), .IN4(n472), .QN(n475) );
  AND2X1 U500 ( .IN1(n231), .IN2(n298), .Q(n230) );
  INVX0 U501 ( .IN(n299), .QN(n231) );
  NAND2X0 U502 ( .IN1(a_in[24]), .IN2(n225), .QN(n232) );
  NBUFFX2 U503 ( .IN(n486), .Q(n247) );
  NBUFFX2 U504 ( .IN(n486), .Q(n246) );
  NBUFFX2 U505 ( .IN(n486), .Q(n245) );
  NBUFFX2 U506 ( .IN(n486), .Q(n244) );
  NBUFFX2 U507 ( .IN(n486), .Q(n243) );
  NBUFFX2 U508 ( .IN(n486), .Q(n242) );
  NBUFFX2 U509 ( .IN(n486), .Q(n241) );
  OR4X1 U510 ( .IN1(reg_b[0]), .IN2(reg_b[10]), .IN3(reg_b[11]), .IN4(
        reg_b[12]), .Q(n70) );
  AO221X1 U511 ( .IN1(n215), .IN2(reg_b[29]), .IN3(a_in[29]), .IN4(n212), 
        .IN5(n467), .Q(N55) );
  AO221X1 U512 ( .IN1(n215), .IN2(reg_b[30]), .IN3(a_in[30]), .IN4(n208), 
        .IN5(n475), .Q(N56) );
  AO221X1 U513 ( .IN1(n492), .IN2(n401), .IN3(n260), .IN4(result[16]), .IN5(
        n400), .Q(N42) );
  AO221X1 U514 ( .IN1(n492), .IN2(n390), .IN3(n261), .IN4(result[14]), .IN5(
        n389), .Q(N40) );
  AO221X1 U515 ( .IN1(n492), .IN2(n398), .IN3(n261), .IN4(result[15]), .IN5(
        n397), .Q(N41) );
  AO221X1 U516 ( .IN1(n492), .IN2(n438), .IN3(n258), .IN4(result[24]), .IN5(
        n437), .Q(N50) );
  AO221X1 U517 ( .IN1(n492), .IN2(n422), .IN3(n259), .IN4(result[20]), .IN5(
        n421), .Q(N46) );
  AO22X1 U518 ( .IN1(a_in[4]), .IN2(n117), .IN3(n215), .IN4(n198), .Q(n343) );
  AO221X1 U519 ( .IN1(n492), .IN2(n482), .IN3(n257), .IN4(result[31]), .IN5(
        n481), .Q(N57) );
  AO22X1 U520 ( .IN1(a_in[31]), .IN2(n117), .IN3(n215), .IN4(reg_b[31]), .Q(
        n481) );
  AO221X1 U521 ( .IN1(n492), .IN2(n383), .IN3(n261), .IN4(result[12]), .IN5(
        n382), .Q(N38) );
  AO22X1 U522 ( .IN1(a_in[12]), .IN2(n118), .IN3(n489), .IN4(reg_b[12]), .Q(
        n382) );
  AO221X1 U523 ( .IN1(n492), .IN2(n410), .IN3(n260), .IN4(result[18]), .IN5(
        n409), .Q(N44) );
  AO22X1 U524 ( .IN1(a_in[18]), .IN2(n117), .IN3(n215), .IN4(reg_b[18]), .Q(
        n409) );
  AO221X1 U525 ( .IN1(n492), .IN2(n454), .IN3(n258), .IN4(result[27]), .IN5(
        n453), .Q(N53) );
  AO22X1 U526 ( .IN1(a_in[27]), .IN2(n118), .IN3(n489), .IN4(reg_b[27]), .Q(
        n453) );
  AO221X1 U527 ( .IN1(n492), .IN2(n432), .IN3(n259), .IN4(result[23]), .IN5(
        n431), .Q(N49) );
  AO22X1 U528 ( .IN1(a_in[23]), .IN2(n224), .IN3(n489), .IN4(reg_b[23]), .Q(
        n431) );
  AO221X1 U529 ( .IN1(n492), .IN2(n371), .IN3(n262), .IN4(result[10]), .IN5(
        n370), .Q(N36) );
  AO22X1 U530 ( .IN1(a_in[10]), .IN2(n118), .IN3(n215), .IN4(reg_b[10]), .Q(
        n370) );
  AO221X1 U531 ( .IN1(n492), .IN2(n426), .IN3(n259), .IN4(result[21]), .IN5(
        n425), .Q(N47) );
  AO22X1 U532 ( .IN1(a_in[21]), .IN2(n117), .IN3(n489), .IN4(reg_b[21]), .Q(
        n425) );
  AO221X1 U533 ( .IN1(n492), .IN2(n418), .IN3(n260), .IN4(result[19]), .IN5(
        n417), .Q(N45) );
  AO22X1 U534 ( .IN1(a_in[19]), .IN2(n117), .IN3(n215), .IN4(reg_b[19]), .Q(
        n417) );
  AO221X1 U535 ( .IN1(n492), .IN2(n484), .IN3(n257), .IN4(result[1]), .IN5(
        n483), .Q(N27) );
  AO22X1 U536 ( .IN1(a_in[1]), .IN2(n118), .IN3(n489), .IN4(n193), .Q(n483) );
  AO221X1 U537 ( .IN1(n492), .IN2(n350), .IN3(n263), .IN4(result[5]), .IN5(
        n349), .Q(N31) );
  AO221X1 U538 ( .IN1(n492), .IN2(n460), .IN3(n257), .IN4(result[28]), .IN5(
        n459), .Q(N54) );
  AO22X1 U539 ( .IN1(a_in[28]), .IN2(n224), .IN3(n489), .IN4(reg_b[28]), .Q(
        n459) );
  AO221X1 U540 ( .IN1(n492), .IN2(n444), .IN3(n258), .IN4(result[25]), .IN5(
        n443), .Q(N51) );
  AO22X1 U541 ( .IN1(a_in[25]), .IN2(n117), .IN3(n489), .IN4(reg_b[25]), .Q(
        n443) );
  AO221X1 U542 ( .IN1(n492), .IN2(n361), .IN3(n262), .IN4(result[8]), .IN5(
        n360), .Q(N34) );
  AO22X1 U543 ( .IN1(a_in[8]), .IN2(n118), .IN3(n489), .IN4(n73), .Q(n360) );
  AO221X1 U544 ( .IN1(n492), .IN2(n405), .IN3(n260), .IN4(result[17]), .IN5(
        n404), .Q(N43) );
  AO22X1 U545 ( .IN1(a_in[17]), .IN2(n118), .IN3(n215), .IN4(reg_b[17]), .Q(
        n404) );
  AO221X1 U546 ( .IN1(n492), .IN2(n379), .IN3(n262), .IN4(result[11]), .IN5(
        n378), .Q(N37) );
  AO22X1 U547 ( .IN1(a_in[11]), .IN2(n117), .IN3(n489), .IN4(reg_b[11]), .Q(
        n378) );
  AO22X1 U548 ( .IN1(a_in[15]), .IN2(n224), .IN3(n215), .IN4(reg_b[15]), .Q(
        n397) );
  AO22X1 U549 ( .IN1(a_in[14]), .IN2(n118), .IN3(n489), .IN4(reg_b[14]), .Q(
        n389) );
  AO22X1 U550 ( .IN1(a_in[16]), .IN2(n224), .IN3(n489), .IN4(reg_b[16]), .Q(
        n400) );
  AO221X1 U551 ( .IN1(n492), .IN2(n449), .IN3(n258), .IN4(result[26]), .IN5(
        n448), .Q(N52) );
  AO22X1 U552 ( .IN1(a_in[26]), .IN2(n224), .IN3(n489), .IN4(reg_b[26]), .Q(
        n448) );
  AO221X1 U553 ( .IN1(n492), .IN2(n429), .IN3(n259), .IN4(result[22]), .IN5(
        n428), .Q(N48) );
  AO22X1 U554 ( .IN1(a_in[22]), .IN2(n118), .IN3(n489), .IN4(reg_b[22]), .Q(
        n428) );
  NOR2X0 U555 ( .IN1(n329), .IN2(n216), .QN(n333) );
  AO222X1 U556 ( .IN1(b_in[4]), .IN2(n249), .IN3(n246), .IN4(n198), .IN5(n237), 
        .IN6(result[4]), .Q(N70) );
  AO221X1 U557 ( .IN1(n492), .IN2(n344), .IN3(n263), .IN4(result[4]), .IN5(
        n343), .Q(N30) );
  NBUFFX2 U558 ( .IN(n486), .Q(n248) );
  AO221X1 U559 ( .IN1(n492), .IN2(n339), .IN3(n257), .IN4(result[3]), .IN5(
        n338), .Q(N29) );
  AO22X1 U560 ( .IN1(a_in[3]), .IN2(n118), .IN3(n489), .IN4(n89), .Q(n338) );
  AO22X1 U561 ( .IN1(a_in[5]), .IN2(n117), .IN3(n489), .IN4(n74), .Q(n349) );
  NOR2X0 U562 ( .IN1(n226), .IN2(n331), .QN(n332) );
  AO222X1 U563 ( .IN1(b_in[0]), .IN2(n253), .IN3(n245), .IN4(reg_b[0]), .IN5(
        n239), .IN6(result[0]), .Q(N66) );
  INVX8 U564 ( .IN(n341), .QN(n282) );
  OAI22X2 U565 ( .IN1(n193), .IN2(n202), .IN3(n97), .IN4(n283), .QN(n324) );
  NAND2X4 U566 ( .IN1(n286), .IN2(n373), .QN(n287) );
  NOR2X4 U567 ( .IN1(n126), .IN2(n303), .QN(n305) );
  NOR2X4 U568 ( .IN1(n305), .IN2(n304), .QN(n306) );
  NAND2X4 U569 ( .IN1(n306), .IN2(n433), .QN(n439) );
  NOR2X4 U570 ( .IN1(n442), .IN2(n307), .QN(n309) );
  NOR2X4 U571 ( .IN1(n309), .IN2(n308), .QN(n310) );
  NAND2X4 U572 ( .IN1(n310), .IN2(n445), .QN(n450) );
  NOR2X4 U573 ( .IN1(n452), .IN2(n311), .QN(n313) );
  NOR2X4 U574 ( .IN1(n313), .IN2(n312), .QN(n314) );
  NAND2X4 U575 ( .IN1(n314), .IN2(n455), .QN(n462) );
  NOR2X4 U576 ( .IN1(n462), .IN2(n315), .QN(n316) );
  NOR2X4 U577 ( .IN1(n316), .IN2(n317), .QN(n320) );
  NAND2X4 U578 ( .IN1(n320), .IN2(n319), .QN(n323) );
endmodule

