module ram_addr_cntr (
        input clk_2,
        input reset_n,
        input ram_ena
        );

endmodule
