module shift_reg (
        input clk_50,
        input reset_n,
        input data_ena,
        input serial_data,
        output [7:0] parallel_data
        );

endmodule
