
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75,
         N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ps;

  AO22X2 U3 ( .IN1(n521), .IN2(gcd_ps[1]), .IN3(n14), .IN4(n15), .Q(n71) );
  NAND2X4 U4 ( .IN1(n16), .IN2(reset_n), .QN(n14) );
  OAI22X2 U5 ( .IN1(n13), .IN2(n15), .IN3(n521), .IN4(n17), .QN(n72) );
  OA21X2 U6 ( .IN1(gcd_ps[1]), .IN2(gcd_ps[0]), .IN3(reset_n), .Q(n17) );
  AO221X2 U9 ( .IN1(start), .IN2(n13), .IN3(n18), .IN4(n520), .IN5(n19), .Q(
        n15) );
  NAND2X4 U10 ( .IN1(reset_n), .IN2(n20), .QN(n19) );
  NAND2X4 U11 ( .IN1(gcd_ps[1]), .IN2(n13), .QN(n20) );
  OR4X4 U118 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n66) );
  OR4X4 U119 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n65) );
  OR4X4 U120 ( .IN1(reg_b[31]), .IN2(reg_b[3]), .IN3(reg_b[4]), .IN4(reg_b[5]), 
        .Q(n64) );
  OR4X4 U121 ( .IN1(reg_b[6]), .IN2(reg_b[7]), .IN3(reg_b[8]), .IN4(reg_b[9]), 
        .Q(n63) );
  OR4X4 U124 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(
        reg_b[16]), .Q(n69) );
  OR4X4 U125 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(
        reg_b[1]), .Q(n68) );
  OR4X4 U126 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n67) );
  DFFARX2 \gcd_ps_reg[0]  ( .D(n72), .CLK(clk), .RSTB(reset_n), .Q(gcd_ps[0]), 
        .QN(n13) );
  DFFARX2 \gcd_ps_reg[1]  ( .D(n71), .CLK(clk), .RSTB(reset_n), .Q(gcd_ps[1]), 
        .QN(n12) );
  DFFX2 \reg_a_reg[1]  ( .D(N27), .CLK(clk), .Q(result[1]) );
  DFFX2 \reg_b_reg[1]  ( .D(N67), .CLK(clk), .Q(reg_b[1]) );
  DFFX2 \reg_a_reg[31]  ( .D(N57), .CLK(clk), .Q(result[31]) );
  DFFX2 \reg_b_reg[31]  ( .D(N97), .CLK(clk), .Q(reg_b[31]) );
  DFFX2 \reg_b_reg[30]  ( .D(N96), .CLK(clk), .Q(reg_b[30]) );
  DFFX2 \reg_a_reg[30]  ( .D(N56), .CLK(clk), .Q(result[30]) );
  DFFX2 \reg_b_reg[29]  ( .D(N95), .CLK(clk), .Q(reg_b[29]) );
  DFFX2 \reg_a_reg[29]  ( .D(N55), .CLK(clk), .Q(result[29]) );
  DFFX2 \reg_b_reg[28]  ( .D(N94), .CLK(clk), .Q(reg_b[28]) );
  DFFX2 \reg_a_reg[28]  ( .D(N54), .CLK(clk), .Q(result[28]) );
  DFFX2 \reg_b_reg[27]  ( .D(N93), .CLK(clk), .Q(reg_b[27]) );
  DFFX2 \reg_a_reg[27]  ( .D(N53), .CLK(clk), .Q(result[27]) );
  DFFX2 \reg_b_reg[26]  ( .D(N92), .CLK(clk), .Q(reg_b[26]) );
  DFFX2 \reg_a_reg[26]  ( .D(N52), .CLK(clk), .Q(result[26]) );
  DFFX2 \reg_b_reg[25]  ( .D(N91), .CLK(clk), .Q(reg_b[25]) );
  DFFX2 \reg_a_reg[25]  ( .D(N51), .CLK(clk), .Q(result[25]) );
  DFFX2 \reg_b_reg[24]  ( .D(N90), .CLK(clk), .Q(reg_b[24]) );
  DFFX2 \reg_a_reg[24]  ( .D(N50), .CLK(clk), .Q(result[24]) );
  DFFX2 \reg_b_reg[23]  ( .D(N89), .CLK(clk), .Q(reg_b[23]) );
  DFFX2 \reg_a_reg[23]  ( .D(N49), .CLK(clk), .Q(result[23]) );
  DFFX2 \reg_b_reg[22]  ( .D(N88), .CLK(clk), .Q(reg_b[22]) );
  DFFX2 \reg_a_reg[22]  ( .D(N48), .CLK(clk), .Q(result[22]) );
  DFFX2 \reg_b_reg[21]  ( .D(N87), .CLK(clk), .Q(reg_b[21]) );
  DFFX2 \reg_a_reg[21]  ( .D(N47), .CLK(clk), .Q(result[21]) );
  DFFX2 \reg_a_reg[20]  ( .D(N46), .CLK(clk), .Q(result[20]) );
  DFFX2 \reg_b_reg[19]  ( .D(N85), .CLK(clk), .Q(reg_b[19]) );
  DFFX2 \reg_a_reg[19]  ( .D(N45), .CLK(clk), .Q(result[19]) );
  DFFX2 \reg_b_reg[18]  ( .D(N84), .CLK(clk), .Q(reg_b[18]) );
  DFFX2 \reg_a_reg[18]  ( .D(N44), .CLK(clk), .Q(result[18]) );
  DFFX2 \reg_b_reg[17]  ( .D(N83), .CLK(clk), .Q(reg_b[17]) );
  DFFX2 \reg_a_reg[17]  ( .D(N43), .CLK(clk), .Q(result[17]) );
  DFFX2 \reg_b_reg[16]  ( .D(N82), .CLK(clk), .Q(reg_b[16]) );
  DFFX2 \reg_a_reg[16]  ( .D(N42), .CLK(clk), .Q(result[16]) );
  DFFX2 \reg_b_reg[15]  ( .D(N81), .CLK(clk), .Q(reg_b[15]) );
  DFFX2 \reg_b_reg[14]  ( .D(N80), .CLK(clk), .Q(reg_b[14]) );
  DFFX2 \reg_a_reg[14]  ( .D(N40), .CLK(clk), .Q(result[14]) );
  DFFX2 \reg_b_reg[13]  ( .D(N79), .CLK(clk), .Q(reg_b[13]) );
  DFFX2 \reg_a_reg[13]  ( .D(N39), .CLK(clk), .Q(result[13]) );
  DFFX2 \reg_b_reg[12]  ( .D(N78), .CLK(clk), .Q(reg_b[12]) );
  DFFX2 \reg_a_reg[12]  ( .D(N38), .CLK(clk), .Q(result[12]) );
  DFFX2 \reg_b_reg[11]  ( .D(N77), .CLK(clk), .Q(reg_b[11]) );
  DFFX2 \reg_a_reg[11]  ( .D(N37), .CLK(clk), .Q(result[11]) );
  DFFX2 \reg_b_reg[10]  ( .D(N76), .CLK(clk), .Q(reg_b[10]) );
  DFFX2 \reg_a_reg[10]  ( .D(N36), .CLK(clk), .Q(result[10]) );
  DFFX2 \reg_b_reg[9]  ( .D(N75), .CLK(clk), .Q(reg_b[9]) );
  DFFX2 \reg_a_reg[9]  ( .D(N35), .CLK(clk), .Q(result[9]) );
  DFFX2 \reg_b_reg[8]  ( .D(N74), .CLK(clk), .Q(reg_b[8]) );
  DFFX2 \reg_a_reg[8]  ( .D(N34), .CLK(clk), .Q(result[8]) );
  DFFX2 \reg_b_reg[7]  ( .D(N73), .CLK(clk), .Q(reg_b[7]) );
  DFFX2 \reg_a_reg[7]  ( .D(N33), .CLK(clk), .Q(result[7]) );
  DFFX2 \reg_b_reg[6]  ( .D(N72), .CLK(clk), .Q(reg_b[6]) );
  DFFX2 \reg_a_reg[6]  ( .D(N32), .CLK(clk), .Q(result[6]) );
  DFFX2 \reg_b_reg[5]  ( .D(N71), .CLK(clk), .Q(reg_b[5]) );
  DFFX2 \reg_a_reg[5]  ( .D(N31), .CLK(clk), .Q(result[5]) );
  DFFX2 \reg_b_reg[4]  ( .D(N70), .CLK(clk), .Q(reg_b[4]) );
  DFFX2 \reg_a_reg[4]  ( .D(N30), .CLK(clk), .Q(result[4]) );
  DFFX2 \reg_b_reg[3]  ( .D(N69), .CLK(clk), .Q(reg_b[3]) );
  DFFX2 \reg_a_reg[3]  ( .D(N29), .CLK(clk), .Q(result[3]) );
  DFFX2 \reg_b_reg[2]  ( .D(N68), .CLK(clk), .Q(reg_b[2]) );
  DFFX2 \reg_a_reg[2]  ( .D(N28), .CLK(clk), .Q(result[2]) );
  DFFX1 \reg_b_reg[0]  ( .D(N66), .CLK(clk), .Q(reg_b[0]) );
  DFFX1 \reg_a_reg[0]  ( .D(N26), .CLK(clk), .Q(result[0]), .QN(n92) );
  DFFX1 \reg_b_reg[20]  ( .D(N86), .CLK(clk), .Q(reg_b[20]), .QN(n77) );
  DFFX1 \reg_a_reg[15]  ( .D(N41), .CLK(clk), .Q(result[15]) );
  INVX1 U135 ( .IN(n98), .QN(n73) );
  INVX2 U136 ( .IN(n96), .QN(n98) );
  INVX8 U137 ( .IN(n96), .QN(n74) );
  INVX8 U138 ( .IN(n74), .QN(n75) );
  OAI22X1 U139 ( .IN1(n76), .IN2(n94), .IN3(n302), .IN4(n77), .QN(n423) );
  INVX32 U140 ( .IN(a_in[20]), .QN(n76) );
  NAND2X2 U141 ( .IN1(n290), .IN2(n293), .QN(n302) );
  NBUFFX2 U142 ( .IN(n517), .Q(n142) );
  INVX8 U143 ( .IN(n94), .QN(n95) );
  INVX1 U144 ( .IN(n98), .QN(n78) );
  INVX2 U145 ( .IN(n138), .QN(n79) );
  NBUFFX2 U146 ( .IN(n517), .Q(n138) );
  INVX8 U147 ( .IN(n82), .QN(n94) );
  NAND2X4 U148 ( .IN1(n512), .IN2(n291), .QN(n496) );
  AND2X2 U149 ( .IN1(n482), .IN2(n483), .Q(n80) );
  OR2X1 U150 ( .IN1(reg_b[28]), .IN2(n144), .Q(n483) );
  INVX4 U151 ( .IN(n85), .QN(n81) );
  INVX8 U152 ( .IN(n84), .QN(n85) );
  OR2X1 U153 ( .IN1(n368), .IN2(n367), .Q(n369) );
  INVX2 U154 ( .IN(n501), .QN(n491) );
  INVX16 U155 ( .IN(n494), .QN(n519) );
  NOR2X4 U156 ( .IN1(n512), .IN2(n293), .QN(n82) );
  NBUFFX16 U157 ( .IN(n517), .Q(n137) );
  INVX4 U158 ( .IN(n302), .QN(n83) );
  INVX8 U159 ( .IN(n302), .QN(n84) );
  INVX8 U160 ( .IN(n302), .QN(n515) );
  NAND2X0 U161 ( .IN1(n519), .IN2(n371), .QN(n86) );
  NAND2X0 U162 ( .IN1(n139), .IN2(result[13]), .QN(n87) );
  INVX2 U163 ( .IN(n370), .QN(n88) );
  NAND3X0 U164 ( .IN1(n86), .IN2(n87), .IN3(n88), .QN(N39) );
  NBUFFX16 U165 ( .IN(n517), .Q(n139) );
  NAND2X0 U166 ( .IN1(n519), .IN2(n330), .QN(n89) );
  NAND2X0 U167 ( .IN1(n141), .IN2(result[7]), .QN(n90) );
  INVX2 U168 ( .IN(n329), .QN(n91) );
  NAND3X0 U169 ( .IN1(n89), .IN2(n90), .IN3(n91), .QN(N33) );
  NBUFFX16 U170 ( .IN(n517), .Q(n141) );
  INVX0 U171 ( .IN(n92), .QN(n93) );
  NOR2X0 U172 ( .IN1(n287), .IN2(n494), .QN(n288) );
  OAI22X1 U173 ( .IN1(n487), .IN2(n496), .IN3(n486), .IN4(n494), .QN(n488) );
  OAI22X1 U174 ( .IN1(n497), .IN2(n496), .IN3(n495), .IN4(n494), .QN(n498) );
  INVX16 U175 ( .IN(n94), .QN(n96) );
  INVX16 U176 ( .IN(n94), .QN(n97) );
  INVX4 U177 ( .IN(n425), .QN(n237) );
  DELLN1X2 U178 ( .IN(n511), .Q(n114) );
  DELLN1X2 U179 ( .IN(n511), .Q(n113) );
  AND2X1 U180 ( .IN1(n381), .IN2(n380), .Q(n384) );
  NAND2X0 U181 ( .IN1(n519), .IN2(n345), .QN(n99) );
  NAND2X0 U182 ( .IN1(n140), .IN2(result[9]), .QN(n100) );
  INVX2 U183 ( .IN(n344), .QN(n101) );
  NAND3X0 U184 ( .IN1(n99), .IN2(n100), .IN3(n101), .QN(N35) );
  NBUFFX16 U185 ( .IN(n517), .Q(n140) );
  NOR2X4 U186 ( .IN1(n217), .IN2(n105), .QN(n102) );
  OR2X2 U187 ( .IN1(n102), .IN2(n103), .Q(n233) );
  AND2X1 U188 ( .IN1(n104), .IN2(n229), .Q(n103) );
  INVX0 U189 ( .IN(n231), .QN(n104) );
  OR2X2 U190 ( .IN1(n413), .IN2(n231), .Q(n105) );
  NAND2X0 U191 ( .IN1(a_in[24]), .IN2(n75), .QN(n106) );
  NAND2X1 U192 ( .IN1(n81), .IN2(reg_b[24]), .QN(n107) );
  NAND2X2 U193 ( .IN1(n106), .IN2(n107), .QN(n451) );
  NBUFFX2 U194 ( .IN(n512), .Q(n123) );
  NBUFFX2 U195 ( .IN(n512), .Q(n122) );
  NBUFFX2 U196 ( .IN(n512), .Q(n121) );
  NBUFFX2 U197 ( .IN(n512), .Q(n120) );
  NBUFFX2 U198 ( .IN(n512), .Q(n119) );
  NBUFFX2 U199 ( .IN(n512), .Q(n118) );
  NBUFFX2 U200 ( .IN(n512), .Q(n117) );
  NBUFFX2 U201 ( .IN(n512), .Q(n124) );
  OR4X1 U202 ( .IN1(reg_b[0]), .IN2(reg_b[10]), .IN3(reg_b[11]), .IN4(
        reg_b[12]), .Q(n70) );
  AO221X1 U203 ( .IN1(n84), .IN2(reg_b[29]), .IN3(a_in[29]), .IN4(n78), .IN5(
        n488), .Q(N55) );
  AO221X1 U204 ( .IN1(n81), .IN2(reg_b[30]), .IN3(a_in[30]), .IN4(n73), .IN5(
        n498), .Q(N56) );
  AO221X1 U205 ( .IN1(n519), .IN2(n393), .IN3(n138), .IN4(result[16]), .IN5(
        n392), .Q(N42) );
  AO221X1 U206 ( .IN1(n519), .IN2(n378), .IN3(n139), .IN4(result[14]), .IN5(
        n377), .Q(N40) );
  AO221X1 U207 ( .IN1(n519), .IN2(n387), .IN3(n139), .IN4(result[15]), .IN5(
        n386), .Q(N41) );
  AO221X1 U208 ( .IN1(n519), .IN2(n452), .IN3(n136), .IN4(result[24]), .IN5(
        n451), .Q(N50) );
  AO221X1 U209 ( .IN1(n519), .IN2(n424), .IN3(n137), .IN4(result[20]), .IN5(
        n423), .Q(N46) );
  AO22X1 U210 ( .IN1(a_in[4]), .IN2(n95), .IN3(n84), .IN4(reg_b[4]), .Q(n310)
         );
  AO221X1 U211 ( .IN1(n519), .IN2(n507), .IN3(n135), .IN4(result[31]), .IN5(
        n506), .Q(N57) );
  AO22X1 U212 ( .IN1(a_in[31]), .IN2(n96), .IN3(n84), .IN4(reg_b[31]), .Q(n506) );
  AO221X1 U213 ( .IN1(n519), .IN2(n366), .IN3(n139), .IN4(result[12]), .IN5(
        n365), .Q(N38) );
  AO22X1 U214 ( .IN1(a_in[12]), .IN2(n95), .IN3(n83), .IN4(reg_b[12]), .Q(n365) );
  AO221X1 U215 ( .IN1(n519), .IN2(n408), .IN3(n138), .IN4(result[18]), .IN5(
        n407), .Q(N44) );
  AO22X1 U216 ( .IN1(a_in[18]), .IN2(n96), .IN3(n84), .IN4(reg_b[18]), .Q(n407) );
  AO221X1 U217 ( .IN1(n519), .IN2(n473), .IN3(n136), .IN4(result[27]), .IN5(
        n472), .Q(N53) );
  AO22X1 U218 ( .IN1(a_in[27]), .IN2(n97), .IN3(n515), .IN4(reg_b[27]), .Q(
        n472) );
  AO221X1 U219 ( .IN1(n519), .IN2(n445), .IN3(n137), .IN4(result[23]), .IN5(
        n444), .Q(N49) );
  AO22X1 U220 ( .IN1(a_in[23]), .IN2(n96), .IN3(n515), .IN4(reg_b[23]), .Q(
        n444) );
  AO221X1 U221 ( .IN1(n519), .IN2(n351), .IN3(n140), .IN4(result[10]), .IN5(
        n350), .Q(N36) );
  AO22X1 U222 ( .IN1(a_in[10]), .IN2(n96), .IN3(n84), .IN4(reg_b[10]), .Q(n350) );
  AO221X1 U223 ( .IN1(n519), .IN2(n325), .IN3(n141), .IN4(result[6]), .IN5(
        n324), .Q(N32) );
  AO22X1 U224 ( .IN1(a_in[6]), .IN2(n95), .IN3(n84), .IN4(reg_b[6]), .Q(n324)
         );
  AO221X1 U225 ( .IN1(n519), .IN2(n431), .IN3(n137), .IN4(result[21]), .IN5(
        n430), .Q(N47) );
  AO22X1 U226 ( .IN1(a_in[21]), .IN2(n96), .IN3(n515), .IN4(reg_b[21]), .Q(
        n430) );
  AO221X1 U227 ( .IN1(n519), .IN2(n417), .IN3(n138), .IN4(result[19]), .IN5(
        n416), .Q(N45) );
  AO22X1 U228 ( .IN1(a_in[19]), .IN2(n95), .IN3(n84), .IN4(reg_b[19]), .Q(n416) );
  AO221X1 U229 ( .IN1(n519), .IN2(n510), .IN3(n135), .IN4(result[1]), .IN5(
        n509), .Q(N27) );
  AO22X1 U230 ( .IN1(a_in[1]), .IN2(n95), .IN3(n83), .IN4(reg_b[1]), .Q(n509)
         );
  AO221X1 U231 ( .IN1(n519), .IN2(n319), .IN3(n141), .IN4(result[5]), .IN5(
        n318), .Q(N31) );
  AO221X1 U232 ( .IN1(n519), .IN2(n518), .IN3(n135), .IN4(n93), .IN5(n516), 
        .Q(N26) );
  AO221X1 U233 ( .IN1(n519), .IN2(n480), .IN3(n135), .IN4(result[28]), .IN5(
        n479), .Q(N54) );
  AO22X1 U234 ( .IN1(a_in[28]), .IN2(n97), .IN3(n515), .IN4(reg_b[28]), .Q(
        n479) );
  AO221X1 U235 ( .IN1(n519), .IN2(n459), .IN3(n136), .IN4(result[25]), .IN5(
        n458), .Q(N51) );
  AO22X1 U236 ( .IN1(a_in[25]), .IN2(n97), .IN3(n515), .IN4(reg_b[25]), .Q(
        n458) );
  AO221X1 U237 ( .IN1(n519), .IN2(n337), .IN3(n140), .IN4(result[8]), .IN5(
        n336), .Q(N34) );
  AO22X1 U238 ( .IN1(a_in[8]), .IN2(n96), .IN3(n83), .IN4(reg_b[8]), .Q(n336)
         );
  AO221X1 U239 ( .IN1(n519), .IN2(n401), .IN3(n138), .IN4(result[17]), .IN5(
        n400), .Q(N43) );
  AO22X1 U240 ( .IN1(a_in[17]), .IN2(n97), .IN3(n84), .IN4(reg_b[17]), .Q(n400) );
  AO221X1 U241 ( .IN1(n519), .IN2(n360), .IN3(n140), .IN4(result[11]), .IN5(
        n359), .Q(N37) );
  AO22X1 U242 ( .IN1(a_in[11]), .IN2(n97), .IN3(n515), .IN4(reg_b[11]), .Q(
        n359) );
  AO22X1 U243 ( .IN1(a_in[13]), .IN2(n75), .IN3(n84), .IN4(reg_b[13]), .Q(n370) );
  AO22X1 U244 ( .IN1(a_in[15]), .IN2(n96), .IN3(n83), .IN4(reg_b[15]), .Q(n386) );
  AO22X1 U245 ( .IN1(a_in[14]), .IN2(n97), .IN3(n83), .IN4(reg_b[14]), .Q(n377) );
  AO22X1 U246 ( .IN1(a_in[16]), .IN2(n95), .IN3(n83), .IN4(reg_b[16]), .Q(n392) );
  INVX4 U247 ( .IN(result[4]), .QN(n186) );
  OAI21X1 U248 ( .IN1(result[4]), .IN2(n200), .IN3(n305), .QN(n315) );
  INVX4 U249 ( .IN(n514), .QN(n508) );
  AO221X1 U250 ( .IN1(n519), .IN2(n466), .IN3(n136), .IN4(result[26]), .IN5(
        n465), .Q(N52) );
  AO221X1 U251 ( .IN1(n204), .IN2(n315), .IN3(reg_b[6]), .IN4(n203), .IN5(n322), .Q(n205) );
  AO22X1 U252 ( .IN1(a_in[26]), .IN2(n97), .IN3(n515), .IN4(reg_b[26]), .Q(
        n465) );
  AO221X1 U253 ( .IN1(n519), .IN2(n438), .IN3(n137), .IN4(result[22]), .IN5(
        n437), .Q(N48) );
  AO22X1 U254 ( .IN1(a_in[22]), .IN2(n97), .IN3(n515), .IN4(reg_b[22]), .Q(
        n437) );
  NOR2X0 U255 ( .IN1(n292), .IN2(n85), .QN(n296) );
  AO222X1 U256 ( .IN1(b_in[4]), .IN2(n126), .IN3(n122), .IN4(reg_b[4]), .IN5(
        n115), .IN6(result[4]), .Q(N70) );
  AO221X1 U257 ( .IN1(n519), .IN2(n311), .IN3(n141), .IN4(result[4]), .IN5(
        n310), .Q(N30) );
  OR2X2 U258 ( .IN1(result[0]), .IN2(n195), .Q(n514) );
  INVX2 U259 ( .IN(reg_b[0]), .QN(n195) );
  NBUFFX2 U260 ( .IN(n512), .Q(n125) );
  AO22X1 U261 ( .IN1(a_in[9]), .IN2(n75), .IN3(n84), .IN4(reg_b[9]), .Q(n344)
         );
  AO22X1 U262 ( .IN1(a_in[7]), .IN2(n75), .IN3(n83), .IN4(reg_b[7]), .Q(n329)
         );
  AO221X1 U263 ( .IN1(n519), .IN2(n304), .IN3(n142), .IN4(result[3]), .IN5(
        n303), .Q(N29) );
  AO22X1 U264 ( .IN1(a_in[3]), .IN2(n97), .IN3(n515), .IN4(reg_b[3]), .Q(n303)
         );
  INVX4 U265 ( .IN(n439), .QN(n246) );
  INVX4 U266 ( .IN(n453), .QN(n255) );
  AO22X1 U267 ( .IN1(a_in[5]), .IN2(n97), .IN3(n515), .IN4(reg_b[5]), .Q(n318)
         );
  OR2X2 U268 ( .IN1(n116), .IN2(n126), .Q(n290) );
  NBUFFX2 U269 ( .IN(n511), .Q(n116) );
  OR3X2 U270 ( .IN1(n379), .IN2(n210), .IN3(n368), .Q(n394) );
  INVX4 U271 ( .IN(n380), .QN(n368) );
  NOR2X0 U272 ( .IN1(n98), .IN2(n294), .QN(n295) );
  AO222X1 U273 ( .IN1(b_in[0]), .IN2(n134), .IN3(n121), .IN4(reg_b[0]), .IN5(
        n108), .IN6(n93), .Q(N66) );
  AO22X1 U274 ( .IN1(a_in[0]), .IN2(n95), .IN3(n83), .IN4(reg_b[0]), .Q(n516)
         );
  OR2X2 U275 ( .IN1(n291), .IN2(n290), .Q(n494) );
  IBUFFX4 U276 ( .IN(n439), .QN(n442) );
  IBUFFX4 U277 ( .IN(n425), .QN(n428) );
  IBUFFX4 U278 ( .IN(n467), .QN(n470) );
  IBUFFX8 U279 ( .IN(n353), .QN(n327) );
  AND2X4 U280 ( .IN1(n354), .IN2(n353), .Q(n357) );
  AND2X4 U281 ( .IN1(n339), .IN2(n353), .Q(n342) );
  NBUFFX32 U282 ( .IN(n511), .Q(n108) );
  NBUFFX32 U283 ( .IN(n511), .Q(n109) );
  NBUFFX32 U284 ( .IN(n511), .Q(n110) );
  NBUFFX32 U285 ( .IN(n511), .Q(n111) );
  NBUFFX32 U286 ( .IN(n511), .Q(n112) );
  NBUFFX32 U287 ( .IN(n511), .Q(n115) );
  NBUFFX32 U288 ( .IN(n513), .Q(n126) );
  NBUFFX32 U289 ( .IN(n513), .Q(n127) );
  NBUFFX32 U290 ( .IN(n513), .Q(n128) );
  NBUFFX32 U291 ( .IN(n513), .Q(n129) );
  NBUFFX32 U292 ( .IN(n513), .Q(n130) );
  NBUFFX32 U293 ( .IN(n513), .Q(n131) );
  NBUFFX32 U294 ( .IN(n513), .Q(n132) );
  NBUFFX32 U295 ( .IN(n513), .Q(n133) );
  NBUFFX32 U296 ( .IN(n513), .Q(n134) );
  NBUFFX32 U297 ( .IN(n517), .Q(n135) );
  NBUFFX32 U298 ( .IN(n517), .Q(n136) );
  INVX8 U299 ( .IN(gcd_ps[0]), .QN(n143) );
  INVX8 U300 ( .IN(n12), .QN(n277) );
  OR2X4 U301 ( .IN1(n143), .IN2(n277), .Q(n16) );
  INVX16 U302 ( .IN(result[2]), .QN(n285) );
  INVX8 U303 ( .IN(result[28]), .QN(n144) );
  INVX16 U304 ( .IN(n483), .QN(n146) );
  INVX8 U305 ( .IN(result[30]), .QN(n497) );
  OR2X4 U306 ( .IN1(reg_b[30]), .IN2(n497), .Q(n499) );
  INVX8 U307 ( .IN(result[29]), .QN(n487) );
  OR2X4 U308 ( .IN1(reg_b[29]), .IN2(n487), .Q(n489) );
  NAND2X4 U309 ( .IN1(n499), .IN2(n489), .QN(n145) );
  NOR2X4 U310 ( .IN1(n146), .IN2(n145), .QN(n150) );
  INVX8 U311 ( .IN(reg_b[29]), .QN(n147) );
  OR2X4 U312 ( .IN1(result[29]), .IN2(n147), .Q(n481) );
  INVX8 U313 ( .IN(n481), .QN(n490) );
  INVX8 U314 ( .IN(result[31]), .QN(n273) );
  INVX8 U315 ( .IN(reg_b[30]), .QN(n148) );
  OR2X4 U316 ( .IN1(result[30]), .IN2(n148), .Q(n500) );
  INVX8 U317 ( .IN(n500), .QN(n149) );
  AO221X2 U318 ( .IN1(n490), .IN2(n499), .IN3(reg_b[31]), .IN4(n273), .IN5(
        n149), .Q(n270) );
  NOR2X4 U319 ( .IN1(n150), .IN2(n270), .QN(n272) );
  INVX8 U320 ( .IN(reg_b[18]), .QN(n152) );
  INVX8 U321 ( .IN(reg_b[17]), .QN(n151) );
  OR2X4 U322 ( .IN1(result[17]), .IN2(n151), .Q(n402) );
  OAI21X2 U323 ( .IN1(result[18]), .IN2(n152), .IN3(n402), .QN(n413) );
  INVX8 U324 ( .IN(result[13]), .QN(n153) );
  OR2X4 U325 ( .IN1(reg_b[13]), .IN2(n153), .Q(n373) );
  INVX8 U326 ( .IN(n373), .QN(n155) );
  INVX8 U327 ( .IN(result[12]), .QN(n176) );
  OR2X4 U328 ( .IN1(reg_b[12]), .IN2(n176), .Q(n154) );
  INVX8 U329 ( .IN(n154), .QN(n367) );
  OR2X4 U330 ( .IN1(n155), .IN2(n367), .Q(n379) );
  INVX8 U331 ( .IN(result[15]), .QN(n156) );
  OR2X4 U332 ( .IN1(reg_b[15]), .IN2(n156), .Q(n388) );
  INVX8 U333 ( .IN(n388), .QN(n159) );
  INVX8 U334 ( .IN(result[14]), .QN(n157) );
  OR2X4 U335 ( .IN1(reg_b[14]), .IN2(n157), .Q(n382) );
  INVX8 U336 ( .IN(n382), .QN(n158) );
  OR2X4 U337 ( .IN1(n159), .IN2(n158), .Q(n210) );
  INVX8 U338 ( .IN(reg_b[11]), .QN(n160) );
  OR2X4 U339 ( .IN1(result[11]), .IN2(n160), .Q(n161) );
  INVX8 U340 ( .IN(n161), .QN(n363) );
  INVX8 U341 ( .IN(result[11]), .QN(n162) );
  OR2X4 U342 ( .IN1(reg_b[11]), .IN2(n162), .Q(n361) );
  INVX8 U343 ( .IN(n361), .QN(n164) );
  INVX8 U344 ( .IN(result[10]), .QN(n173) );
  OR2X4 U345 ( .IN1(reg_b[10]), .IN2(n173), .Q(n355) );
  INVX8 U346 ( .IN(n355), .QN(n163) );
  OR2X4 U347 ( .IN1(n164), .IN2(n163), .Q(n184) );
  INVX8 U348 ( .IN(n184), .QN(n175) );
  INVX8 U349 ( .IN(result[9]), .QN(n165) );
  OR2X4 U350 ( .IN1(reg_b[9]), .IN2(n165), .Q(n346) );
  INVX8 U351 ( .IN(n346), .QN(n168) );
  INVX8 U352 ( .IN(result[8]), .QN(n166) );
  OR2X4 U353 ( .IN1(reg_b[8]), .IN2(n166), .Q(n340) );
  INVX8 U354 ( .IN(n340), .QN(n167) );
  OR2X4 U355 ( .IN1(n168), .IN2(n167), .Q(n183) );
  INVX8 U356 ( .IN(n183), .QN(n174) );
  INVX8 U357 ( .IN(reg_b[8]), .QN(n170) );
  INVX8 U358 ( .IN(reg_b[7]), .QN(n169) );
  OR2X4 U359 ( .IN1(result[7]), .IN2(n169), .Q(n331) );
  OAI21X2 U360 ( .IN1(result[8]), .IN2(n170), .IN3(n331), .QN(n341) );
  INVX8 U361 ( .IN(reg_b[9]), .QN(n171) );
  OR2X4 U362 ( .IN1(result[9]), .IN2(n171), .Q(n172) );
  INVX8 U363 ( .IN(n172), .QN(n348) );
  AO221X2 U364 ( .IN1(n174), .IN2(n341), .IN3(reg_b[10]), .IN4(n173), .IN5(
        n348), .Q(n356) );
  NAND2X4 U365 ( .IN1(n175), .IN2(n356), .QN(n178) );
  NAND2X4 U366 ( .IN1(reg_b[12]), .IN2(n176), .QN(n177) );
  NAND2X4 U367 ( .IN1(n178), .IN2(n177), .QN(n179) );
  NOR2X4 U368 ( .IN1(n363), .IN2(n179), .QN(n209) );
  INVX8 U369 ( .IN(result[7]), .QN(n180) );
  OR2X4 U370 ( .IN1(reg_b[7]), .IN2(n180), .Q(n332) );
  INVX8 U371 ( .IN(n332), .QN(n182) );
  INVX8 U372 ( .IN(result[6]), .QN(n203) );
  OR2X4 U373 ( .IN1(reg_b[6]), .IN2(n203), .Q(n181) );
  INVX8 U374 ( .IN(n181), .QN(n326) );
  OR2X4 U375 ( .IN1(n182), .IN2(n326), .Q(n338) );
  OR2X4 U376 ( .IN1(n338), .IN2(n183), .Q(n352) );
  NOR2X4 U377 ( .IN1(n352), .IN2(n184), .QN(n207) );
  INVX8 U378 ( .IN(result[5]), .QN(n185) );
  OR2X4 U379 ( .IN1(reg_b[5]), .IN2(n185), .Q(n320) );
  INVX8 U380 ( .IN(n320), .QN(n188) );
  OR2X4 U381 ( .IN1(reg_b[4]), .IN2(n186), .Q(n314) );
  INVX8 U382 ( .IN(n314), .QN(n187) );
  OR2X4 U383 ( .IN1(n188), .IN2(n187), .Q(n189) );
  INVX8 U384 ( .IN(n189), .QN(n204) );
  INVX8 U385 ( .IN(result[3]), .QN(n190) );
  OR2X4 U386 ( .IN1(reg_b[3]), .IN2(n190), .Q(n306) );
  INVX8 U387 ( .IN(n306), .QN(n193) );
  INVX8 U388 ( .IN(result[2]), .QN(n191) );
  OR2X4 U389 ( .IN1(reg_b[2]), .IN2(n191), .Q(n192) );
  INVX8 U390 ( .IN(n192), .QN(n299) );
  OR2X4 U391 ( .IN1(n193), .IN2(n299), .Q(n194) );
  INVX8 U392 ( .IN(n194), .QN(n313) );
  AND2X2 U393 ( .IN1(n204), .IN2(n313), .Q(n206) );
  INVX8 U394 ( .IN(reg_b[2]), .QN(n198) );
  INVX8 U395 ( .IN(result[1]), .QN(n197) );
  AND2X2 U396 ( .IN1(reg_b[1]), .IN2(n197), .Q(n196) );
  OAI22X2 U397 ( .IN1(reg_b[1]), .IN2(n197), .IN3(n508), .IN4(n196), .QN(n286)
         );
  OAI21X2 U398 ( .IN1(result[2]), .IN2(n198), .IN3(n286), .QN(n312) );
  INVX8 U399 ( .IN(reg_b[4]), .QN(n200) );
  INVX8 U400 ( .IN(reg_b[3]), .QN(n199) );
  OR2X4 U401 ( .IN1(result[3]), .IN2(n199), .Q(n305) );
  INVX8 U402 ( .IN(reg_b[5]), .QN(n201) );
  OR2X4 U403 ( .IN1(result[5]), .IN2(n201), .Q(n202) );
  INVX8 U404 ( .IN(n202), .QN(n322) );
  AO21X2 U405 ( .IN1(n206), .IN2(n312), .IN3(n205), .Q(n353) );
  NAND2X4 U406 ( .IN1(n207), .IN2(n353), .QN(n208) );
  NAND2X4 U407 ( .IN1(n208), .IN2(n209), .QN(n380) );
  INVX8 U408 ( .IN(n210), .QN(n215) );
  INVX8 U409 ( .IN(reg_b[14]), .QN(n212) );
  INVX8 U410 ( .IN(reg_b[13]), .QN(n211) );
  OR2X4 U411 ( .IN1(result[13]), .IN2(n211), .Q(n372) );
  OAI21X2 U412 ( .IN1(result[14]), .IN2(n212), .IN3(n372), .QN(n383) );
  INVX8 U413 ( .IN(result[16]), .QN(n223) );
  INVX8 U414 ( .IN(reg_b[15]), .QN(n213) );
  OR2X4 U415 ( .IN1(result[15]), .IN2(n213), .Q(n214) );
  INVX8 U416 ( .IN(n214), .QN(n390) );
  AO221X2 U417 ( .IN1(n215), .IN2(n383), .IN3(reg_b[16]), .IN4(n223), .IN5(
        n390), .Q(n395) );
  INVX16 U418 ( .IN(n395), .QN(n216) );
  NAND2X4 U419 ( .IN1(n394), .IN2(n216), .QN(n217) );
  INVX8 U420 ( .IN(result[19]), .QN(n218) );
  OR2X4 U421 ( .IN1(reg_b[19]), .IN2(n218), .Q(n419) );
  INVX16 U422 ( .IN(n419), .QN(n221) );
  INVX8 U423 ( .IN(result[18]), .QN(n219) );
  OR2X4 U424 ( .IN1(reg_b[18]), .IN2(n219), .Q(n412) );
  INVX16 U425 ( .IN(n412), .QN(n220) );
  NOR2X4 U426 ( .IN1(n221), .IN2(n220), .QN(n228) );
  INVX8 U427 ( .IN(result[17]), .QN(n222) );
  OR2X4 U428 ( .IN1(reg_b[17]), .IN2(n222), .Q(n403) );
  INVX8 U429 ( .IN(n403), .QN(n225) );
  OR2X4 U430 ( .IN1(reg_b[16]), .IN2(n223), .Q(n224) );
  INVX8 U431 ( .IN(n224), .QN(n398) );
  OR2X4 U432 ( .IN1(n225), .IN2(n398), .Q(n409) );
  INVX16 U433 ( .IN(n413), .QN(n226) );
  NAND2X4 U434 ( .IN1(n409), .IN2(n226), .QN(n227) );
  NAND2X4 U435 ( .IN1(n228), .IN2(n227), .QN(n229) );
  INVX16 U436 ( .IN(reg_b[20]), .QN(n230) );
  NOR2X4 U437 ( .IN1(result[20]), .IN2(n230), .QN(n231) );
  INVX8 U438 ( .IN(reg_b[19]), .QN(n232) );
  OR2X4 U439 ( .IN1(result[19]), .IN2(n232), .Q(n418) );
  NAND2X4 U440 ( .IN1(n233), .IN2(n418), .QN(n425) );
  INVX8 U441 ( .IN(result[20]), .QN(n234) );
  OR2X4 U442 ( .IN1(reg_b[20]), .IN2(n234), .Q(n426) );
  INVX8 U443 ( .IN(result[21]), .QN(n235) );
  OR2X4 U444 ( .IN1(reg_b[21]), .IN2(n235), .Q(n433) );
  NAND2X4 U445 ( .IN1(n426), .IN2(n433), .QN(n236) );
  NOR2X4 U446 ( .IN1(n237), .IN2(n236), .QN(n240) );
  INVX16 U447 ( .IN(reg_b[22]), .QN(n238) );
  NOR2X4 U448 ( .IN1(result[22]), .IN2(n238), .QN(n239) );
  NOR2X4 U449 ( .IN1(n240), .IN2(n239), .QN(n242) );
  INVX8 U450 ( .IN(reg_b[21]), .QN(n241) );
  OR2X4 U451 ( .IN1(result[21]), .IN2(n241), .Q(n432) );
  NAND2X4 U452 ( .IN1(n242), .IN2(n432), .QN(n439) );
  INVX8 U453 ( .IN(result[22]), .QN(n243) );
  OR2X4 U454 ( .IN1(reg_b[22]), .IN2(n243), .Q(n440) );
  INVX8 U455 ( .IN(result[23]), .QN(n244) );
  OR2X4 U456 ( .IN1(reg_b[23]), .IN2(n244), .Q(n447) );
  NAND2X4 U457 ( .IN1(n440), .IN2(n447), .QN(n245) );
  NOR2X4 U458 ( .IN1(n246), .IN2(n245), .QN(n249) );
  INVX16 U459 ( .IN(reg_b[24]), .QN(n247) );
  NOR2X4 U460 ( .IN1(result[24]), .IN2(n247), .QN(n248) );
  NOR2X4 U461 ( .IN1(n249), .IN2(n248), .QN(n251) );
  INVX8 U462 ( .IN(reg_b[23]), .QN(n250) );
  OR2X4 U463 ( .IN1(result[23]), .IN2(n250), .Q(n446) );
  NAND2X4 U464 ( .IN1(n251), .IN2(n446), .QN(n453) );
  INVX8 U465 ( .IN(result[24]), .QN(n252) );
  OR2X4 U466 ( .IN1(reg_b[24]), .IN2(n252), .Q(n454) );
  INVX8 U467 ( .IN(result[25]), .QN(n253) );
  OR2X4 U468 ( .IN1(reg_b[25]), .IN2(n253), .Q(n461) );
  NAND2X4 U469 ( .IN1(n454), .IN2(n461), .QN(n254) );
  NOR2X4 U470 ( .IN1(n255), .IN2(n254), .QN(n258) );
  INVX16 U471 ( .IN(reg_b[26]), .QN(n256) );
  NOR2X4 U472 ( .IN1(result[26]), .IN2(n256), .QN(n257) );
  NOR2X4 U473 ( .IN1(n258), .IN2(n257), .QN(n260) );
  INVX8 U474 ( .IN(reg_b[25]), .QN(n259) );
  OR2X4 U475 ( .IN1(result[25]), .IN2(n259), .Q(n460) );
  NAND2X4 U476 ( .IN1(n260), .IN2(n460), .QN(n467) );
  INVX16 U477 ( .IN(n467), .QN(n264) );
  INVX8 U478 ( .IN(result[26]), .QN(n261) );
  OR2X4 U479 ( .IN1(reg_b[26]), .IN2(n261), .Q(n468) );
  INVX8 U480 ( .IN(result[27]), .QN(n262) );
  OR2X4 U481 ( .IN1(reg_b[27]), .IN2(n262), .Q(n475) );
  NAND2X4 U482 ( .IN1(n468), .IN2(n475), .QN(n263) );
  NOR2X4 U483 ( .IN1(n264), .IN2(n263), .QN(n267) );
  INVX16 U484 ( .IN(reg_b[28]), .QN(n265) );
  NOR2X4 U485 ( .IN1(result[28]), .IN2(n265), .QN(n266) );
  NOR2X4 U486 ( .IN1(n267), .IN2(n266), .QN(n269) );
  INVX8 U487 ( .IN(reg_b[27]), .QN(n268) );
  OR2X4 U488 ( .IN1(result[27]), .IN2(n268), .Q(n474) );
  NAND2X4 U489 ( .IN1(n269), .IN2(n474), .QN(n482) );
  NOR2X4 U490 ( .IN1(n482), .IN2(n270), .QN(n271) );
  NOR2X4 U491 ( .IN1(n272), .IN2(n271), .QN(n276) );
  OR2X4 U492 ( .IN1(reg_b[31]), .IN2(n273), .Q(n502) );
  INVX16 U493 ( .IN(n502), .QN(n274) );
  NOR2X4 U494 ( .IN1(n16), .IN2(n274), .QN(n275) );
  NAND2X4 U495 ( .IN1(n276), .IN2(n275), .QN(n284) );
  INVX8 U496 ( .IN(n284), .QN(n511) );
  INVX8 U497 ( .IN(start), .QN(n279) );
  INVX8 U498 ( .IN(n13), .QN(n278) );
  OR3X4 U499 ( .IN1(n279), .IN2(n278), .IN3(n277), .Q(n280) );
  INVX8 U500 ( .IN(n280), .QN(n513) );
  OR4X2 U501 ( .IN1(n64), .IN2(n63), .IN3(n66), .IN4(n65), .Q(n282) );
  OR4X2 U502 ( .IN1(n68), .IN2(n67), .IN3(n70), .IN4(n69), .Q(n281) );
  OR2X4 U503 ( .IN1(n282), .IN2(n281), .Q(n283) );
  INVX8 U504 ( .IN(n283), .QN(n18) );
  OAI21X2 U505 ( .IN1(n16), .IN2(n18), .IN3(n284), .QN(n293) );
  NOR2X4 U506 ( .IN1(n285), .IN2(n79), .QN(n289) );
  XOR3X2 U507 ( .IN1(result[2]), .IN2(n286), .IN3(reg_b[2]), .Q(n287) );
  INVX8 U508 ( .IN(n293), .QN(n291) );
  NOR2X4 U509 ( .IN1(n289), .IN2(n288), .QN(n298) );
  INVX16 U510 ( .IN(reg_b[2]), .QN(n292) );
  INVX8 U511 ( .IN(n290), .QN(n512) );
  INVX16 U512 ( .IN(a_in[2]), .QN(n294) );
  NOR2X4 U513 ( .IN1(n296), .IN2(n295), .QN(n297) );
  NAND2X4 U514 ( .IN1(n298), .IN2(n297), .QN(N28) );
  AO222X2 U515 ( .IN1(b_in[2]), .IN2(n126), .IN3(n123), .IN4(reg_b[2]), .IN5(
        n115), .IN6(result[2]), .Q(N68) );
  INVX8 U516 ( .IN(n312), .QN(n300) );
  OR2X4 U517 ( .IN1(n300), .IN2(n299), .Q(n301) );
  INVX8 U518 ( .IN(n301), .QN(n307) );
  XOR3X2 U519 ( .IN1(result[3]), .IN2(reg_b[3]), .IN3(n307), .Q(n304) );
  INVX8 U520 ( .IN(n496), .QN(n517) );
  AO222X2 U521 ( .IN1(b_in[3]), .IN2(n126), .IN3(n122), .IN4(reg_b[3]), .IN5(
        n115), .IN6(result[3]), .Q(N69) );
  INVX8 U522 ( .IN(n305), .QN(n308) );
  OA21X2 U523 ( .IN1(n308), .IN2(n307), .IN3(n306), .Q(n309) );
  XOR3X2 U524 ( .IN1(result[4]), .IN2(reg_b[4]), .IN3(n309), .Q(n311) );
  AND2X2 U525 ( .IN1(n313), .IN2(n312), .Q(n316) );
  OAI21X2 U526 ( .IN1(n316), .IN2(n315), .IN3(n314), .QN(n317) );
  INVX8 U527 ( .IN(n317), .QN(n321) );
  XOR3X2 U528 ( .IN1(result[5]), .IN2(reg_b[5]), .IN3(n321), .Q(n319) );
  AO222X2 U529 ( .IN1(b_in[5]), .IN2(n127), .IN3(n121), .IN4(reg_b[5]), .IN5(
        n115), .IN6(result[5]), .Q(N71) );
  OA21X2 U530 ( .IN1(n322), .IN2(n321), .IN3(n320), .Q(n323) );
  XOR3X2 U531 ( .IN1(reg_b[6]), .IN2(result[6]), .IN3(n323), .Q(n325) );
  AO222X2 U532 ( .IN1(b_in[6]), .IN2(n127), .IN3(n120), .IN4(reg_b[6]), .IN5(
        n114), .IN6(result[6]), .Q(N72) );
  OR2X4 U533 ( .IN1(n327), .IN2(n326), .Q(n328) );
  INVX8 U534 ( .IN(n328), .QN(n333) );
  XOR3X2 U535 ( .IN1(result[7]), .IN2(reg_b[7]), .IN3(n333), .Q(n330) );
  AO222X2 U536 ( .IN1(b_in[7]), .IN2(n127), .IN3(n119), .IN4(reg_b[7]), .IN5(
        n114), .IN6(result[7]), .Q(N73) );
  INVX8 U537 ( .IN(n331), .QN(n334) );
  OA21X2 U538 ( .IN1(n334), .IN2(n333), .IN3(n332), .Q(n335) );
  XOR3X2 U539 ( .IN1(result[8]), .IN2(reg_b[8]), .IN3(n335), .Q(n337) );
  AO222X2 U540 ( .IN1(b_in[8]), .IN2(n127), .IN3(n118), .IN4(reg_b[8]), .IN5(
        n114), .IN6(result[8]), .Q(N74) );
  INVX8 U541 ( .IN(n338), .QN(n339) );
  OAI21X2 U542 ( .IN1(n342), .IN2(n341), .IN3(n340), .QN(n343) );
  INVX8 U543 ( .IN(n343), .QN(n347) );
  XOR3X2 U544 ( .IN1(result[9]), .IN2(reg_b[9]), .IN3(n347), .Q(n345) );
  AO222X2 U545 ( .IN1(b_in[9]), .IN2(n128), .IN3(n117), .IN4(reg_b[9]), .IN5(
        n114), .IN6(result[9]), .Q(N75) );
  OA21X2 U546 ( .IN1(n348), .IN2(n347), .IN3(n346), .Q(n349) );
  XOR3X2 U547 ( .IN1(result[10]), .IN2(reg_b[10]), .IN3(n349), .Q(n351) );
  AO222X2 U548 ( .IN1(b_in[10]), .IN2(n128), .IN3(n124), .IN4(reg_b[10]), 
        .IN5(n113), .IN6(result[10]), .Q(N76) );
  INVX8 U549 ( .IN(n352), .QN(n354) );
  OAI21X2 U550 ( .IN1(n357), .IN2(n356), .IN3(n355), .QN(n358) );
  INVX8 U551 ( .IN(n358), .QN(n362) );
  XOR3X2 U552 ( .IN1(result[11]), .IN2(reg_b[11]), .IN3(n362), .Q(n360) );
  AO222X2 U553 ( .IN1(b_in[11]), .IN2(n128), .IN3(n123), .IN4(reg_b[11]), 
        .IN5(n113), .IN6(result[11]), .Q(N77) );
  OA21X2 U554 ( .IN1(n363), .IN2(n362), .IN3(n361), .Q(n364) );
  XOR3X2 U555 ( .IN1(reg_b[12]), .IN2(result[12]), .IN3(n364), .Q(n366) );
  AO222X2 U556 ( .IN1(b_in[12]), .IN2(n128), .IN3(n122), .IN4(reg_b[12]), 
        .IN5(n113), .IN6(result[12]), .Q(N78) );
  INVX8 U557 ( .IN(n369), .QN(n374) );
  XOR3X2 U558 ( .IN1(result[13]), .IN2(reg_b[13]), .IN3(n374), .Q(n371) );
  AO222X2 U559 ( .IN1(b_in[13]), .IN2(n129), .IN3(n121), .IN4(reg_b[13]), 
        .IN5(n113), .IN6(result[13]), .Q(N79) );
  INVX8 U560 ( .IN(n372), .QN(n375) );
  OA21X2 U561 ( .IN1(n375), .IN2(n374), .IN3(n373), .Q(n376) );
  XOR3X2 U562 ( .IN1(result[14]), .IN2(reg_b[14]), .IN3(n376), .Q(n378) );
  AO222X2 U563 ( .IN1(b_in[14]), .IN2(n129), .IN3(n120), .IN4(reg_b[14]), 
        .IN5(n112), .IN6(result[14]), .Q(N80) );
  INVX8 U564 ( .IN(n379), .QN(n381) );
  OAI21X2 U565 ( .IN1(n384), .IN2(n383), .IN3(n382), .QN(n385) );
  INVX8 U566 ( .IN(n385), .QN(n389) );
  XOR3X2 U567 ( .IN1(result[15]), .IN2(reg_b[15]), .IN3(n389), .Q(n387) );
  AO222X2 U568 ( .IN1(b_in[15]), .IN2(n129), .IN3(n119), .IN4(reg_b[15]), 
        .IN5(n112), .IN6(result[15]), .Q(N81) );
  OA21X2 U569 ( .IN1(n390), .IN2(n389), .IN3(n388), .Q(n391) );
  XOR3X2 U570 ( .IN1(result[16]), .IN2(reg_b[16]), .IN3(n391), .Q(n393) );
  AO222X2 U571 ( .IN1(b_in[16]), .IN2(n129), .IN3(n118), .IN4(reg_b[16]), 
        .IN5(n112), .IN6(result[16]), .Q(N82) );
  INVX8 U572 ( .IN(n394), .QN(n396) );
  OR2X4 U573 ( .IN1(n396), .IN2(n395), .Q(n410) );
  INVX8 U574 ( .IN(n410), .QN(n397) );
  OR2X4 U575 ( .IN1(n398), .IN2(n397), .Q(n399) );
  INVX8 U576 ( .IN(n399), .QN(n404) );
  XOR3X2 U577 ( .IN1(result[17]), .IN2(reg_b[17]), .IN3(n404), .Q(n401) );
  AO222X2 U578 ( .IN1(b_in[17]), .IN2(n130), .IN3(n117), .IN4(reg_b[17]), 
        .IN5(n112), .IN6(result[17]), .Q(N83) );
  INVX8 U579 ( .IN(n402), .QN(n405) );
  OA21X2 U580 ( .IN1(n405), .IN2(n404), .IN3(n403), .Q(n406) );
  XOR3X2 U581 ( .IN1(reg_b[18]), .IN2(result[18]), .IN3(n406), .Q(n408) );
  AO222X2 U582 ( .IN1(b_in[18]), .IN2(n130), .IN3(n118), .IN4(reg_b[18]), 
        .IN5(n111), .IN6(result[18]), .Q(N84) );
  INVX8 U583 ( .IN(n409), .QN(n411) );
  AND2X2 U584 ( .IN1(n411), .IN2(n410), .Q(n414) );
  OAI21X2 U585 ( .IN1(n414), .IN2(n413), .IN3(n412), .QN(n415) );
  INVX8 U586 ( .IN(n415), .QN(n420) );
  XOR3X2 U587 ( .IN1(result[19]), .IN2(reg_b[19]), .IN3(n420), .Q(n417) );
  AO222X2 U588 ( .IN1(b_in[19]), .IN2(n130), .IN3(n117), .IN4(reg_b[19]), 
        .IN5(n111), .IN6(result[19]), .Q(N85) );
  INVX8 U589 ( .IN(n418), .QN(n421) );
  OA21X2 U590 ( .IN1(n421), .IN2(n420), .IN3(n419), .Q(n422) );
  XOR3X2 U591 ( .IN1(reg_b[20]), .IN2(result[20]), .IN3(n422), .Q(n424) );
  AO222X2 U592 ( .IN1(b_in[20]), .IN2(n130), .IN3(n124), .IN4(reg_b[20]), 
        .IN5(n111), .IN6(result[20]), .Q(N86) );
  INVX8 U593 ( .IN(n426), .QN(n427) );
  OR2X4 U594 ( .IN1(n428), .IN2(n427), .Q(n429) );
  INVX8 U595 ( .IN(n429), .QN(n434) );
  XOR3X2 U596 ( .IN1(result[21]), .IN2(reg_b[21]), .IN3(n434), .Q(n431) );
  AO222X2 U597 ( .IN1(b_in[21]), .IN2(n131), .IN3(n125), .IN4(reg_b[21]), 
        .IN5(n111), .IN6(result[21]), .Q(N87) );
  INVX8 U598 ( .IN(n432), .QN(n435) );
  OA21X2 U599 ( .IN1(n435), .IN2(n434), .IN3(n433), .Q(n436) );
  XOR3X2 U600 ( .IN1(reg_b[22]), .IN2(result[22]), .IN3(n436), .Q(n438) );
  AO222X2 U601 ( .IN1(b_in[22]), .IN2(n131), .IN3(n122), .IN4(reg_b[22]), 
        .IN5(n110), .IN6(result[22]), .Q(N88) );
  INVX8 U602 ( .IN(n440), .QN(n441) );
  OR2X4 U603 ( .IN1(n442), .IN2(n441), .Q(n443) );
  INVX8 U604 ( .IN(n443), .QN(n448) );
  XOR3X2 U605 ( .IN1(result[23]), .IN2(reg_b[23]), .IN3(n448), .Q(n445) );
  AO222X2 U606 ( .IN1(b_in[23]), .IN2(n131), .IN3(n121), .IN4(reg_b[23]), 
        .IN5(n110), .IN6(result[23]), .Q(N89) );
  INVX8 U607 ( .IN(n446), .QN(n449) );
  OA21X2 U608 ( .IN1(n449), .IN2(n448), .IN3(n447), .Q(n450) );
  XOR3X2 U609 ( .IN1(reg_b[24]), .IN2(result[24]), .IN3(n450), .Q(n452) );
  AO222X2 U610 ( .IN1(b_in[24]), .IN2(n131), .IN3(n120), .IN4(reg_b[24]), 
        .IN5(n110), .IN6(result[24]), .Q(N90) );
  INVX8 U611 ( .IN(n453), .QN(n456) );
  INVX8 U612 ( .IN(n454), .QN(n455) );
  OR2X4 U613 ( .IN1(n456), .IN2(n455), .Q(n457) );
  INVX8 U614 ( .IN(n457), .QN(n462) );
  XOR3X2 U615 ( .IN1(result[25]), .IN2(reg_b[25]), .IN3(n462), .Q(n459) );
  AO222X2 U616 ( .IN1(b_in[25]), .IN2(n132), .IN3(n119), .IN4(reg_b[25]), 
        .IN5(n110), .IN6(result[25]), .Q(N91) );
  INVX8 U617 ( .IN(n460), .QN(n463) );
  OA21X2 U618 ( .IN1(n463), .IN2(n462), .IN3(n461), .Q(n464) );
  XOR3X2 U619 ( .IN1(reg_b[26]), .IN2(result[26]), .IN3(n464), .Q(n466) );
  AO222X2 U620 ( .IN1(b_in[26]), .IN2(n132), .IN3(n125), .IN4(reg_b[26]), 
        .IN5(n109), .IN6(result[26]), .Q(N92) );
  INVX8 U621 ( .IN(n468), .QN(n469) );
  OR2X4 U622 ( .IN1(n470), .IN2(n469), .Q(n471) );
  INVX8 U623 ( .IN(n471), .QN(n476) );
  XOR3X2 U624 ( .IN1(result[27]), .IN2(reg_b[27]), .IN3(n476), .Q(n473) );
  AO222X2 U625 ( .IN1(b_in[27]), .IN2(n132), .IN3(n125), .IN4(reg_b[27]), 
        .IN5(n109), .IN6(result[27]), .Q(N93) );
  INVX8 U626 ( .IN(n474), .QN(n477) );
  OA21X2 U627 ( .IN1(n477), .IN2(n476), .IN3(n475), .Q(n478) );
  XOR3X2 U628 ( .IN1(reg_b[28]), .IN2(result[28]), .IN3(n478), .Q(n480) );
  AO222X2 U629 ( .IN1(b_in[28]), .IN2(n132), .IN3(n125), .IN4(reg_b[28]), 
        .IN5(n109), .IN6(result[28]), .Q(N94) );
  AND2X2 U630 ( .IN1(n481), .IN2(n489), .Q(n485) );
  XOR2X2 U631 ( .IN1(result[29]), .IN2(reg_b[29]), .Q(n484) );
  MUX21X2 U632 ( .IN1(n485), .IN2(n484), .S(n80), .Q(n486) );
  AO222X2 U633 ( .IN1(b_in[29]), .IN2(n133), .IN3(n123), .IN4(reg_b[29]), 
        .IN5(n109), .IN6(result[29]), .Q(N95) );
  AND2X2 U634 ( .IN1(n500), .IN2(n499), .Q(n493) );
  XOR2X2 U635 ( .IN1(result[30]), .IN2(reg_b[30]), .Q(n492) );
  OAI21X2 U636 ( .IN1(n490), .IN2(n80), .IN3(n489), .QN(n501) );
  MUX21X2 U637 ( .IN1(n493), .IN2(n492), .S(n491), .Q(n495) );
  AO222X2 U638 ( .IN1(b_in[30]), .IN2(n133), .IN3(n124), .IN4(reg_b[30]), 
        .IN5(n108), .IN6(result[30]), .Q(N96) );
  AO222X2 U639 ( .IN1(b_in[31]), .IN2(n133), .IN3(n125), .IN4(reg_b[31]), 
        .IN5(n108), .IN6(result[31]), .Q(N97) );
  INVX8 U640 ( .IN(n499), .QN(n505) );
  AND2X2 U641 ( .IN1(n501), .IN2(n500), .Q(n504) );
  INVX8 U642 ( .IN(n502), .QN(n503) );
  OA21X2 U643 ( .IN1(n505), .IN2(n504), .IN3(n503), .Q(n507) );
  AO222X2 U644 ( .IN1(b_in[1]), .IN2(n133), .IN3(n123), .IN4(reg_b[1]), .IN5(
        n108), .IN6(result[1]), .Q(N67) );
  XOR3X2 U645 ( .IN1(reg_b[1]), .IN2(result[1]), .IN3(n508), .Q(n510) );
  OAI21X2 U646 ( .IN1(reg_b[0]), .IN2(n92), .IN3(n514), .QN(n518) );
  INVX8 U647 ( .IN(n16), .QN(n520) );
  INVX16 U648 ( .IN(n15), .QN(n521) );
  INVX16 U649 ( .IN(n20), .QN(done) );
endmodule

