module ctrl_blk_50(
	input 		a5_or_c3,
	input 		data_ena,
	input 		clk_50,
	input 		reset_n,
	output reg 	wr_fifo);

enum reg {not_detect	= 1'b0,
          detect	= 1'b1,
          detect_xx	= 'x} detect_ps, detect_ns;

enum reg {not_write	= 1'b0,
          write		= 1'b1,
          write_xx	= 'x} write_ps, write_ns;

enum reg [2:0]  {	header	= 3'b000,
          		data_0	= 3'b001,
	  		data_1	= 3'b010,
	  		data_2	= 3'b011,
	  		data_3	= 3'b100,
          		data_type_xx	= 'x} data_type_ps, data_type_ns;

enum reg {check		= 1'b0,
          temp		= 1'b1,
          packet_xx	= 'x} packet_type_ps, packet_type_ns;


wire byte_assembled;
wire [1:0] packet_cntr;

//assignmants
assign byte_assembled = ((detect_ps) & (!data_ena)) ? 1'b1 : 1'b0; 

//************************************************************
//sm #1  Is there data on the serial data line?
//************************************************************
always_ff @(posedge clk_50, negedge reset_n)
    	if (!reset_n) detect_ps <= not_detect;        //after reset, go to state 'not_complete'
    	else          detect_ps <= detect_ns;        //else, go to next state

always_comb begin
    	detect_ns = detect_xx;   //default assignments
         
    	case (detect_ps)
     		not_detect:
      			if (data_ena == 1'b1) 	detect_ns = detect;
      			else               	detect_ns = not_detect;
     		detect:
      			if (data_ena == 1'b1) 	detect_ns = detect;
      			else               	detect_ns = not_detect;
    	endcase
end//always_comb


//************************************************************
//sm #2 packet type
//************************************************************
always_ff @(posedge clk_50, negedge reset_n)
    	if (!reset_n) packet_type_ps <= check;        	
    	else          packet_type_ps <= packet_type_ns;        //else, go to next state

always_comb begin
    	packet_type_ns = packet_xx;   //default assignments
         
    	case (packet_type_ps)
     		check:
			if ((data_type_ps == header) & (a5_or_c3) & (byte_assembled)) packet_type_ns = temp;
			else packet_type_ns = check;

     		temp:
      			if (data_type_ps != header ) 	packet_type_ns = temp; 
      			else 				packet_type_ns = check; 
    	endcase
end//always_comb



//************************************************************
//sm #3 header or data 
//************************************************************
always_ff @(posedge clk_50, negedge reset_n)
    	if (!reset_n) data_type_ps <= header;        //after reset, go to state 'not_complete'
    	else          data_type_ps <= data_type_ns;        //else, go to next state

always_comb begin
    	data_type_ns = data_type_xx;   //default assignments
         
    	case (data_type_ps)
     		header:
			if ( byte_assembled ) 	data_type_ns = data_0;
			else			data_type_ns = header;	
     		data_0:
      			if ( byte_assembled ) 	data_type_ns = data_1;
      			else 			data_type_ns = data_0; 
     		data_1:
      			if ( byte_assembled ) 	data_type_ns = data_2;
      			else 			data_type_ns = data_1; 
     		data_2:
      			if ( byte_assembled ) 	data_type_ns = data_3;
      			else 			data_type_ns = data_2; 
     		data_3:
      			if ( byte_assembled ) 	data_type_ns = header;
      			else 			data_type_ns = data_3; 
    	endcase
end//always_comb


//************************************************************
//sm #4 write state
//************************************************************
always_ff @(posedge clk_50, negedge reset_n)
    	if (!reset_n) write_ps <= not_write;        	
    	else          write_ps <= write_ns;        //else, go to next state

always_comb begin
    	write_ns = write_xx;   //default assignments
        wr_fifo = 1'b0;
    	case (write_ps)
     		not_write:
			if  ((data_type_ps != header) & (packet_type_ps == temp) & (byte_assembled)) write_ns = write;
			else write_ns = not_write;

     		write:
			begin
				wr_fifo = 1'b1;
      				write_ns = not_write; 
			end
    	endcase
end//always_comb


endmodule
