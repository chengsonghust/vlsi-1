module accumulator (
        input  data_in,
        input  zero_select,
        input  rd_fifo,
        input  clk_2,
        input  reset_n,
        output [8:0] acc_out
        );

endmodule
